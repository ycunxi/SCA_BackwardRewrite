// Benchmark "CSAMultiplier" written by ABC on Tue Sep 16 13:49:27 2014

module CSAMultiplier ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , b0 ,
    b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 , b9 ,
    b10 , b11 , b12 , b13 , b14 , b15 ,
    z0 , z1 , z2 , z3 , z4 , z5 , z6 , z7 , z8 ,
    z9 , z10 , z11 , z12 , z13 , z14 , z15 , z16 ,
    z17 , z18 , z19 , z20 , z21 , z22 , z23 , z24 ,
    z25 , z26 , z27 , z28 , z29 , z30 , z31   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    b0 , b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 ,
    b9 , b10 , b11 , b12 , b13 , b14 , b15 ;
  output z0 , z1 , z2 , z3 , z4 , z5 , z6 , z7 ,
    z8 , z9 , z10 , z11 , z12 , z13 , z14 , z15 ,
    z16 , z17 , z18 , z19 , z20 , z21 , z22 , z23 ,
    z24 , z25 , z26 , z27 , z28 , z29 , z30 , z31 ;
  wire n65, n66, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2266, n2267, n2268, n2269;
  and2  g0000(.a(b0 ), .b(a0 ), .O(z0 ));
  and2  g0001(.a(b1 ), .b(a0 ), .O(n65));
  and2  g0002(.a(b0 ), .b(a1 ), .O(n66));
  xor2  g0003(.a(n66), .b(n65), .O(z1 ));
  and2  g0004(.a(b2 ), .b(a0 ), .O(n68));
  and2  g0005(.a(n66), .b(n65), .O(n69));
  xor2  g0006(.a(n69), .b(n68), .O(n70));
  and2  g0007(.a(b1 ), .b(a1 ), .O(n71));
  and2  g0008(.a(b0 ), .b(a2 ), .O(n72));
  xor2  g0009(.a(n72), .b(n71), .O(n73));
  xor2  g0010(.a(n73), .b(n70), .O(z2 ));
  nand2 g0011(.a(b3 ), .b(a0 ), .O(n75));
  inv1  g0012(.a(n75), .O(n76));
  nand2 g0013(.a(n73), .b(n69), .O(n77));
  nand2 g0014(.a(n69), .b(n68), .O(n78));
  nand2 g0015(.a(n73), .b(n68), .O(n79));
  and2  g0016(.a(n79), .b(n78), .O(n80));
  nand2 g0017(.a(n80), .b(n77), .O(n81));
  xor2  g0018(.a(n81), .b(n76), .O(n82));
  nand2 g0019(.a(b2 ), .b(a1 ), .O(n83));
  and2  g0020(.a(b1 ), .b(a2 ), .O(n84));
  and2  g0021(.a(b0 ), .b(a3 ), .O(n85));
  xor2  g0022(.a(n85), .b(n84), .O(n86));
  xor2  g0023(.a(n86), .b(n83), .O(n87));
  nand2 g0024(.a(n72), .b(n71), .O(n88));
  xor2  g0025(.a(n88), .b(n87), .O(n89));
  xor2  g0026(.a(n89), .b(n82), .O(z3 ));
  nand2 g0027(.a(b4 ), .b(a0 ), .O(n91));
  inv1  g0028(.a(n91), .O(n92));
  nand2 g0029(.a(n89), .b(n81), .O(n93));
  nand2 g0030(.a(n81), .b(n76), .O(n94));
  nand2 g0031(.a(n89), .b(n76), .O(n95));
  and2  g0032(.a(n95), .b(n94), .O(n96));
  nand2 g0033(.a(n96), .b(n93), .O(n97));
  xor2  g0034(.a(n97), .b(n92), .O(n98));
  nand2 g0035(.a(b3 ), .b(a1 ), .O(n99));
  inv1  g0036(.a(n99), .O(n100));
  nand2 g0037(.a(b2 ), .b(a2 ), .O(n101));
  inv1  g0038(.a(n101), .O(n102));
  and2  g0039(.a(b1 ), .b(a3 ), .O(n103));
  and2  g0040(.a(b0 ), .b(a4 ), .O(n104));
  xor2  g0041(.a(n104), .b(n103), .O(n105));
  xor2  g0042(.a(n105), .b(n102), .O(n106));
  and2  g0043(.a(n85), .b(n84), .O(n107));
  xor2  g0044(.a(n107), .b(n106), .O(n108));
  xor2  g0045(.a(n108), .b(n100), .O(n109));
  inv1  g0046(.a(n88), .O(n110));
  nand2 g0047(.a(n110), .b(n86), .O(n111));
  inv1  g0048(.a(n83), .O(n112));
  nand2 g0049(.a(n110), .b(n112), .O(n113));
  nand2 g0050(.a(n86), .b(n112), .O(n114));
  and2  g0051(.a(n114), .b(n113), .O(n115));
  nand2 g0052(.a(n115), .b(n111), .O(n116));
  xor2  g0053(.a(n116), .b(n109), .O(n117));
  xor2  g0054(.a(n117), .b(n98), .O(z4 ));
  nand2 g0055(.a(b5 ), .b(a0 ), .O(n119));
  inv1  g0056(.a(n119), .O(n120));
  nand2 g0057(.a(n117), .b(n97), .O(n121));
  nand2 g0058(.a(n97), .b(n92), .O(n122));
  nand2 g0059(.a(n117), .b(n92), .O(n123));
  and2  g0060(.a(n123), .b(n122), .O(n124));
  nand2 g0061(.a(n124), .b(n121), .O(n125));
  xor2  g0062(.a(n125), .b(n120), .O(n126));
  nand2 g0063(.a(b4 ), .b(a1 ), .O(n127));
  inv1  g0064(.a(n127), .O(n128));
  nand2 g0065(.a(b3 ), .b(a2 ), .O(n129));
  inv1  g0066(.a(n129), .O(n130));
  nand2 g0067(.a(b2 ), .b(a3 ), .O(n131));
  inv1  g0068(.a(n131), .O(n132));
  and2  g0069(.a(b1 ), .b(a4 ), .O(n133));
  and2  g0070(.a(b0 ), .b(a5 ), .O(n134));
  xor2  g0071(.a(n134), .b(n133), .O(n135));
  xor2  g0072(.a(n135), .b(n132), .O(n136));
  and2  g0073(.a(n104), .b(n103), .O(n137));
  xor2  g0074(.a(n137), .b(n136), .O(n138));
  xor2  g0075(.a(n138), .b(n130), .O(n139));
  nand2 g0076(.a(n107), .b(n105), .O(n140));
  nand2 g0077(.a(n107), .b(n102), .O(n141));
  nand2 g0078(.a(n105), .b(n102), .O(n142));
  and2  g0079(.a(n142), .b(n141), .O(n143));
  nand2 g0080(.a(n143), .b(n140), .O(n144));
  xor2  g0081(.a(n144), .b(n139), .O(n145));
  xor2  g0082(.a(n145), .b(n128), .O(n146));
  nand2 g0083(.a(n116), .b(n108), .O(n147));
  nand2 g0084(.a(n116), .b(n100), .O(n148));
  nand2 g0085(.a(n108), .b(n100), .O(n149));
  and2  g0086(.a(n149), .b(n148), .O(n150));
  nand2 g0087(.a(n150), .b(n147), .O(n151));
  xor2  g0088(.a(n151), .b(n146), .O(n152));
  xor2  g0089(.a(n152), .b(n126), .O(z5 ));
  nand2 g0090(.a(b6 ), .b(a0 ), .O(n154));
  inv1  g0091(.a(n154), .O(n155));
  nand2 g0092(.a(n152), .b(n125), .O(n156));
  nand2 g0093(.a(n125), .b(n120), .O(n157));
  nand2 g0094(.a(n152), .b(n120), .O(n158));
  and2  g0095(.a(n158), .b(n157), .O(n159));
  nand2 g0096(.a(n159), .b(n156), .O(n160));
  xor2  g0097(.a(n160), .b(n155), .O(n161));
  nand2 g0098(.a(b5 ), .b(a1 ), .O(n162));
  inv1  g0099(.a(n162), .O(n163));
  nand2 g0100(.a(b4 ), .b(a2 ), .O(n164));
  inv1  g0101(.a(n164), .O(n165));
  nand2 g0102(.a(b3 ), .b(a3 ), .O(n166));
  inv1  g0103(.a(n166), .O(n167));
  nand2 g0104(.a(b2 ), .b(a4 ), .O(n168));
  inv1  g0105(.a(n168), .O(n169));
  and2  g0106(.a(b1 ), .b(a5 ), .O(n170));
  and2  g0107(.a(b0 ), .b(a6 ), .O(n171));
  xor2  g0108(.a(n171), .b(n170), .O(n172));
  xor2  g0109(.a(n172), .b(n169), .O(n173));
  and2  g0110(.a(n134), .b(n133), .O(n174));
  xor2  g0111(.a(n174), .b(n173), .O(n175));
  xor2  g0112(.a(n175), .b(n167), .O(n176));
  nand2 g0113(.a(n137), .b(n135), .O(n177));
  nand2 g0114(.a(n137), .b(n132), .O(n178));
  nand2 g0115(.a(n135), .b(n132), .O(n179));
  and2  g0116(.a(n179), .b(n178), .O(n180));
  nand2 g0117(.a(n180), .b(n177), .O(n181));
  xor2  g0118(.a(n181), .b(n176), .O(n182));
  xor2  g0119(.a(n182), .b(n165), .O(n183));
  nand2 g0120(.a(n144), .b(n138), .O(n184));
  nand2 g0121(.a(n144), .b(n130), .O(n185));
  nand2 g0122(.a(n138), .b(n130), .O(n186));
  and2  g0123(.a(n186), .b(n185), .O(n187));
  nand2 g0124(.a(n187), .b(n184), .O(n188));
  xor2  g0125(.a(n188), .b(n183), .O(n189));
  xor2  g0126(.a(n189), .b(n163), .O(n190));
  nand2 g0127(.a(n151), .b(n145), .O(n191));
  nand2 g0128(.a(n151), .b(n128), .O(n192));
  nand2 g0129(.a(n145), .b(n128), .O(n193));
  and2  g0130(.a(n193), .b(n192), .O(n194));
  nand2 g0131(.a(n194), .b(n191), .O(n195));
  xor2  g0132(.a(n195), .b(n190), .O(n196));
  xor2  g0133(.a(n196), .b(n161), .O(z6 ));
  nand2 g0134(.a(b7 ), .b(a0 ), .O(n198));
  inv1  g0135(.a(n198), .O(n199));
  nand2 g0136(.a(n196), .b(n160), .O(n200));
  nand2 g0137(.a(n160), .b(n155), .O(n201));
  nand2 g0138(.a(n196), .b(n155), .O(n202));
  and2  g0139(.a(n202), .b(n201), .O(n203));
  nand2 g0140(.a(n203), .b(n200), .O(n204));
  xor2  g0141(.a(n204), .b(n199), .O(n205));
  nand2 g0142(.a(b6 ), .b(a1 ), .O(n206));
  nand2 g0143(.a(b5 ), .b(a2 ), .O(n207));
  nand2 g0144(.a(b4 ), .b(a3 ), .O(n208));
  inv1  g0145(.a(n208), .O(n209));
  nand2 g0146(.a(b3 ), .b(a4 ), .O(n210));
  inv1  g0147(.a(n210), .O(n211));
  nand2 g0148(.a(b2 ), .b(a5 ), .O(n212));
  inv1  g0149(.a(n212), .O(n213));
  and2  g0150(.a(b1 ), .b(a6 ), .O(n214));
  and2  g0151(.a(b0 ), .b(a7 ), .O(n215));
  xor2  g0152(.a(n215), .b(n214), .O(n216));
  xor2  g0153(.a(n216), .b(n213), .O(n217));
  and2  g0154(.a(n171), .b(n170), .O(n218));
  xor2  g0155(.a(n218), .b(n217), .O(n219));
  xor2  g0156(.a(n219), .b(n211), .O(n220));
  nand2 g0157(.a(n174), .b(n172), .O(n221));
  nand2 g0158(.a(n174), .b(n169), .O(n222));
  nand2 g0159(.a(n172), .b(n169), .O(n223));
  and2  g0160(.a(n223), .b(n222), .O(n224));
  nand2 g0161(.a(n224), .b(n221), .O(n225));
  xor2  g0162(.a(n225), .b(n220), .O(n226));
  xor2  g0163(.a(n226), .b(n209), .O(n227));
  nand2 g0164(.a(n181), .b(n175), .O(n228));
  nand2 g0165(.a(n181), .b(n167), .O(n229));
  nand2 g0166(.a(n175), .b(n167), .O(n230));
  and2  g0167(.a(n230), .b(n229), .O(n231));
  nand2 g0168(.a(n231), .b(n228), .O(n232));
  xor2  g0169(.a(n232), .b(n227), .O(n233));
  xor2  g0170(.a(n233), .b(n207), .O(n234));
  nand2 g0171(.a(n188), .b(n182), .O(n235));
  nand2 g0172(.a(n188), .b(n165), .O(n236));
  nand2 g0173(.a(n182), .b(n165), .O(n237));
  and2  g0174(.a(n237), .b(n236), .O(n238));
  nand2 g0175(.a(n238), .b(n235), .O(n239));
  xor2  g0176(.a(n239), .b(n234), .O(n240));
  xor2  g0177(.a(n240), .b(n206), .O(n241));
  nand2 g0178(.a(n195), .b(n189), .O(n242));
  nand2 g0179(.a(n195), .b(n163), .O(n243));
  nand2 g0180(.a(n189), .b(n163), .O(n244));
  and2  g0181(.a(n244), .b(n243), .O(n245));
  nand2 g0182(.a(n245), .b(n242), .O(n246));
  xor2  g0183(.a(n246), .b(n241), .O(n247));
  xor2  g0184(.a(n247), .b(n205), .O(z7 ));
  nand2 g0185(.a(b8 ), .b(a0 ), .O(n249));
  inv1  g0186(.a(n249), .O(n250));
  nand2 g0187(.a(n247), .b(n204), .O(n251));
  nand2 g0188(.a(n204), .b(n199), .O(n252));
  nand2 g0189(.a(n247), .b(n199), .O(n253));
  and2  g0190(.a(n253), .b(n252), .O(n254));
  nand2 g0191(.a(n254), .b(n251), .O(n255));
  xor2  g0192(.a(n255), .b(n250), .O(n256));
  nand2 g0193(.a(b7 ), .b(a1 ), .O(n257));
  nand2 g0194(.a(b6 ), .b(a2 ), .O(n258));
  nand2 g0195(.a(b5 ), .b(a3 ), .O(n259));
  inv1  g0196(.a(n259), .O(n260));
  nand2 g0197(.a(b4 ), .b(a4 ), .O(n261));
  inv1  g0198(.a(n261), .O(n262));
  nand2 g0199(.a(b3 ), .b(a5 ), .O(n263));
  inv1  g0200(.a(n263), .O(n264));
  nand2 g0201(.a(b2 ), .b(a6 ), .O(n265));
  inv1  g0202(.a(n265), .O(n266));
  and2  g0203(.a(b1 ), .b(a7 ), .O(n267));
  and2  g0204(.a(b0 ), .b(a8 ), .O(n268));
  xor2  g0205(.a(n268), .b(n267), .O(n269));
  xor2  g0206(.a(n269), .b(n266), .O(n270));
  and2  g0207(.a(n215), .b(n214), .O(n271));
  xor2  g0208(.a(n271), .b(n270), .O(n272));
  xor2  g0209(.a(n272), .b(n264), .O(n273));
  nand2 g0210(.a(n218), .b(n216), .O(n274));
  nand2 g0211(.a(n218), .b(n213), .O(n275));
  nand2 g0212(.a(n216), .b(n213), .O(n276));
  and2  g0213(.a(n276), .b(n275), .O(n277));
  nand2 g0214(.a(n277), .b(n274), .O(n278));
  xor2  g0215(.a(n278), .b(n273), .O(n279));
  xor2  g0216(.a(n279), .b(n262), .O(n280));
  nand2 g0217(.a(n225), .b(n219), .O(n281));
  nand2 g0218(.a(n225), .b(n211), .O(n282));
  nand2 g0219(.a(n219), .b(n211), .O(n283));
  and2  g0220(.a(n283), .b(n282), .O(n284));
  nand2 g0221(.a(n284), .b(n281), .O(n285));
  xor2  g0222(.a(n285), .b(n280), .O(n286));
  xor2  g0223(.a(n286), .b(n260), .O(n287));
  nand2 g0224(.a(n232), .b(n226), .O(n288));
  nand2 g0225(.a(n232), .b(n209), .O(n289));
  nand2 g0226(.a(n226), .b(n209), .O(n290));
  and2  g0227(.a(n290), .b(n289), .O(n291));
  nand2 g0228(.a(n291), .b(n288), .O(n292));
  xor2  g0229(.a(n292), .b(n287), .O(n293));
  xor2  g0230(.a(n293), .b(n258), .O(n294));
  nand2 g0231(.a(n239), .b(n233), .O(n295));
  inv1  g0232(.a(n207), .O(n296));
  nand2 g0233(.a(n239), .b(n296), .O(n297));
  nand2 g0234(.a(n233), .b(n296), .O(n298));
  and2  g0235(.a(n298), .b(n297), .O(n299));
  nand2 g0236(.a(n299), .b(n295), .O(n300));
  xor2  g0237(.a(n300), .b(n294), .O(n301));
  xor2  g0238(.a(n301), .b(n257), .O(n302));
  inv1  g0239(.a(n240), .O(n303));
  nand2 g0240(.a(n246), .b(n303), .O(n304));
  inv1  g0241(.a(n206), .O(n305));
  nand2 g0242(.a(n246), .b(n305), .O(n306));
  nand2 g0243(.a(n303), .b(n305), .O(n307));
  and2  g0244(.a(n307), .b(n306), .O(n308));
  nand2 g0245(.a(n308), .b(n304), .O(n309));
  xor2  g0246(.a(n309), .b(n302), .O(n310));
  xor2  g0247(.a(n310), .b(n256), .O(z8 ));
  nand2 g0248(.a(b9 ), .b(a0 ), .O(n312));
  inv1  g0249(.a(n312), .O(n313));
  nand2 g0250(.a(n310), .b(n255), .O(n314));
  nand2 g0251(.a(n255), .b(n250), .O(n315));
  nand2 g0252(.a(n310), .b(n250), .O(n316));
  and2  g0253(.a(n316), .b(n315), .O(n317));
  nand2 g0254(.a(n317), .b(n314), .O(n318));
  xor2  g0255(.a(n318), .b(n313), .O(n319));
  nand2 g0256(.a(b8 ), .b(a1 ), .O(n320));
  nand2 g0257(.a(b7 ), .b(a2 ), .O(n321));
  nand2 g0258(.a(b6 ), .b(a3 ), .O(n322));
  inv1  g0259(.a(n322), .O(n323));
  nand2 g0260(.a(b5 ), .b(a4 ), .O(n324));
  inv1  g0261(.a(n324), .O(n325));
  nand2 g0262(.a(b4 ), .b(a5 ), .O(n326));
  inv1  g0263(.a(n326), .O(n327));
  nand2 g0264(.a(b3 ), .b(a6 ), .O(n328));
  inv1  g0265(.a(n328), .O(n329));
  nand2 g0266(.a(b2 ), .b(a7 ), .O(n330));
  inv1  g0267(.a(n330), .O(n331));
  and2  g0268(.a(b1 ), .b(a8 ), .O(n332));
  and2  g0269(.a(b0 ), .b(a9 ), .O(n333));
  xor2  g0270(.a(n333), .b(n332), .O(n334));
  xor2  g0271(.a(n334), .b(n331), .O(n335));
  and2  g0272(.a(n268), .b(n267), .O(n336));
  xor2  g0273(.a(n336), .b(n335), .O(n337));
  xor2  g0274(.a(n337), .b(n329), .O(n338));
  nand2 g0275(.a(n271), .b(n269), .O(n339));
  nand2 g0276(.a(n271), .b(n266), .O(n340));
  nand2 g0277(.a(n269), .b(n266), .O(n341));
  and2  g0278(.a(n341), .b(n340), .O(n342));
  nand2 g0279(.a(n342), .b(n339), .O(n343));
  xor2  g0280(.a(n343), .b(n338), .O(n344));
  xor2  g0281(.a(n344), .b(n327), .O(n345));
  nand2 g0282(.a(n278), .b(n272), .O(n346));
  nand2 g0283(.a(n278), .b(n264), .O(n347));
  nand2 g0284(.a(n272), .b(n264), .O(n348));
  and2  g0285(.a(n348), .b(n347), .O(n349));
  nand2 g0286(.a(n349), .b(n346), .O(n350));
  xor2  g0287(.a(n350), .b(n345), .O(n351));
  xor2  g0288(.a(n351), .b(n325), .O(n352));
  nand2 g0289(.a(n285), .b(n279), .O(n353));
  nand2 g0290(.a(n285), .b(n262), .O(n354));
  nand2 g0291(.a(n279), .b(n262), .O(n355));
  and2  g0292(.a(n355), .b(n354), .O(n356));
  nand2 g0293(.a(n356), .b(n353), .O(n357));
  xor2  g0294(.a(n357), .b(n352), .O(n358));
  xor2  g0295(.a(n358), .b(n323), .O(n359));
  nand2 g0296(.a(n292), .b(n286), .O(n360));
  nand2 g0297(.a(n292), .b(n260), .O(n361));
  nand2 g0298(.a(n286), .b(n260), .O(n362));
  and2  g0299(.a(n362), .b(n361), .O(n363));
  nand2 g0300(.a(n363), .b(n360), .O(n364));
  xor2  g0301(.a(n364), .b(n359), .O(n365));
  xor2  g0302(.a(n365), .b(n321), .O(n366));
  nand2 g0303(.a(n300), .b(n293), .O(n367));
  inv1  g0304(.a(n258), .O(n368));
  nand2 g0305(.a(n300), .b(n368), .O(n369));
  nand2 g0306(.a(n293), .b(n368), .O(n370));
  and2  g0307(.a(n370), .b(n369), .O(n371));
  nand2 g0308(.a(n371), .b(n367), .O(n372));
  xor2  g0309(.a(n372), .b(n366), .O(n373));
  xor2  g0310(.a(n373), .b(n320), .O(n374));
  inv1  g0311(.a(n301), .O(n375));
  nand2 g0312(.a(n309), .b(n375), .O(n376));
  inv1  g0313(.a(n257), .O(n377));
  nand2 g0314(.a(n309), .b(n377), .O(n378));
  nand2 g0315(.a(n375), .b(n377), .O(n379));
  and2  g0316(.a(n379), .b(n378), .O(n380));
  nand2 g0317(.a(n380), .b(n376), .O(n381));
  xor2  g0318(.a(n381), .b(n374), .O(n382));
  xor2  g0319(.a(n382), .b(n319), .O(z9 ));
  nand2 g0320(.a(b10 ), .b(a0 ), .O(n384));
  inv1  g0321(.a(n384), .O(n385));
  nand2 g0322(.a(n382), .b(n318), .O(n386));
  nand2 g0323(.a(n318), .b(n313), .O(n387));
  nand2 g0324(.a(n382), .b(n313), .O(n388));
  and2  g0325(.a(n388), .b(n387), .O(n389));
  nand2 g0326(.a(n389), .b(n386), .O(n390));
  xor2  g0327(.a(n390), .b(n385), .O(n391));
  nand2 g0328(.a(b9 ), .b(a1 ), .O(n392));
  inv1  g0329(.a(n392), .O(n393));
  nand2 g0330(.a(b8 ), .b(a2 ), .O(n394));
  inv1  g0331(.a(n394), .O(n395));
  nand2 g0332(.a(b7 ), .b(a3 ), .O(n396));
  inv1  g0333(.a(n396), .O(n397));
  nand2 g0334(.a(b6 ), .b(a4 ), .O(n398));
  inv1  g0335(.a(n398), .O(n399));
  nand2 g0336(.a(b5 ), .b(a5 ), .O(n400));
  inv1  g0337(.a(n400), .O(n401));
  nand2 g0338(.a(b4 ), .b(a6 ), .O(n402));
  inv1  g0339(.a(n402), .O(n403));
  nand2 g0340(.a(b3 ), .b(a7 ), .O(n404));
  inv1  g0341(.a(n404), .O(n405));
  nand2 g0342(.a(b2 ), .b(a8 ), .O(n406));
  inv1  g0343(.a(n406), .O(n407));
  nand2 g0344(.a(b1 ), .b(a9 ), .O(n408));
  nand2 g0345(.a(b0 ), .b(a10 ), .O(n409));
  xor2  g0346(.a(n409), .b(n408), .O(n410));
  xor2  g0347(.a(n410), .b(n407), .O(n411));
  and2  g0348(.a(n333), .b(n332), .O(n412));
  xor2  g0349(.a(n412), .b(n411), .O(n413));
  xor2  g0350(.a(n413), .b(n405), .O(n414));
  nand2 g0351(.a(n336), .b(n334), .O(n415));
  nand2 g0352(.a(n336), .b(n331), .O(n416));
  nand2 g0353(.a(n334), .b(n331), .O(n417));
  and2  g0354(.a(n417), .b(n416), .O(n418));
  nand2 g0355(.a(n418), .b(n415), .O(n419));
  xor2  g0356(.a(n419), .b(n414), .O(n420));
  xor2  g0357(.a(n420), .b(n403), .O(n421));
  nand2 g0358(.a(n343), .b(n337), .O(n422));
  nand2 g0359(.a(n343), .b(n329), .O(n423));
  nand2 g0360(.a(n337), .b(n329), .O(n424));
  and2  g0361(.a(n424), .b(n423), .O(n425));
  nand2 g0362(.a(n425), .b(n422), .O(n426));
  xor2  g0363(.a(n426), .b(n421), .O(n427));
  xor2  g0364(.a(n427), .b(n401), .O(n428));
  nand2 g0365(.a(n350), .b(n344), .O(n429));
  nand2 g0366(.a(n350), .b(n327), .O(n430));
  nand2 g0367(.a(n344), .b(n327), .O(n431));
  and2  g0368(.a(n431), .b(n430), .O(n432));
  nand2 g0369(.a(n432), .b(n429), .O(n433));
  xor2  g0370(.a(n433), .b(n428), .O(n434));
  xor2  g0371(.a(n434), .b(n399), .O(n435));
  nand2 g0372(.a(n357), .b(n351), .O(n436));
  nand2 g0373(.a(n357), .b(n325), .O(n437));
  nand2 g0374(.a(n351), .b(n325), .O(n438));
  and2  g0375(.a(n438), .b(n437), .O(n439));
  nand2 g0376(.a(n439), .b(n436), .O(n440));
  xor2  g0377(.a(n440), .b(n435), .O(n441));
  xor2  g0378(.a(n441), .b(n397), .O(n442));
  nand2 g0379(.a(n364), .b(n358), .O(n443));
  nand2 g0380(.a(n364), .b(n323), .O(n444));
  nand2 g0381(.a(n358), .b(n323), .O(n445));
  and2  g0382(.a(n445), .b(n444), .O(n446));
  nand2 g0383(.a(n446), .b(n443), .O(n447));
  xor2  g0384(.a(n447), .b(n442), .O(n448));
  xor2  g0385(.a(n448), .b(n395), .O(n449));
  nand2 g0386(.a(n372), .b(n365), .O(n450));
  inv1  g0387(.a(n321), .O(n451));
  nand2 g0388(.a(n372), .b(n451), .O(n452));
  nand2 g0389(.a(n365), .b(n451), .O(n453));
  and2  g0390(.a(n453), .b(n452), .O(n454));
  nand2 g0391(.a(n454), .b(n450), .O(n455));
  xor2  g0392(.a(n455), .b(n449), .O(n456));
  xor2  g0393(.a(n456), .b(n393), .O(n457));
  inv1  g0394(.a(n373), .O(n458));
  nand2 g0395(.a(n381), .b(n458), .O(n459));
  inv1  g0396(.a(n320), .O(n460));
  nand2 g0397(.a(n381), .b(n460), .O(n461));
  nand2 g0398(.a(n458), .b(n460), .O(n462));
  and2  g0399(.a(n462), .b(n461), .O(n463));
  nand2 g0400(.a(n463), .b(n459), .O(n464));
  xor2  g0401(.a(n464), .b(n457), .O(n465));
  xor2  g0402(.a(n465), .b(n391), .O(z10 ));
  nand2 g0403(.a(b11 ), .b(a0 ), .O(n467));
  inv1  g0404(.a(n467), .O(n468));
  nand2 g0405(.a(n465), .b(n390), .O(n469));
  nand2 g0406(.a(n390), .b(n385), .O(n470));
  nand2 g0407(.a(n465), .b(n385), .O(n471));
  and2  g0408(.a(n471), .b(n470), .O(n472));
  nand2 g0409(.a(n472), .b(n469), .O(n473));
  xor2  g0410(.a(n473), .b(n468), .O(n474));
  nand2 g0411(.a(b10 ), .b(a1 ), .O(n475));
  inv1  g0412(.a(n475), .O(n476));
  nand2 g0413(.a(b9 ), .b(a2 ), .O(n477));
  inv1  g0414(.a(n477), .O(n478));
  nand2 g0415(.a(b8 ), .b(a3 ), .O(n479));
  inv1  g0416(.a(n479), .O(n480));
  nand2 g0417(.a(b7 ), .b(a4 ), .O(n481));
  inv1  g0418(.a(n481), .O(n482));
  nand2 g0419(.a(b6 ), .b(a5 ), .O(n483));
  inv1  g0420(.a(n483), .O(n484));
  nand2 g0421(.a(b5 ), .b(a6 ), .O(n485));
  inv1  g0422(.a(n485), .O(n486));
  nand2 g0423(.a(b4 ), .b(a7 ), .O(n487));
  inv1  g0424(.a(n487), .O(n488));
  nand2 g0425(.a(b3 ), .b(a8 ), .O(n489));
  inv1  g0426(.a(n489), .O(n490));
  nand2 g0427(.a(b2 ), .b(a9 ), .O(n491));
  inv1  g0428(.a(n491), .O(n492));
  nand2 g0429(.a(b1 ), .b(a10 ), .O(n493));
  nand2 g0430(.a(b0 ), .b(a11 ), .O(n494));
  xor2  g0431(.a(n494), .b(n493), .O(n495));
  xor2  g0432(.a(n495), .b(n492), .O(n496));
  or2   g0433(.a(n409), .b(n408), .O(n497));
  inv1  g0434(.a(n497), .O(n498));
  xor2  g0435(.a(n498), .b(n496), .O(n499));
  xor2  g0436(.a(n499), .b(n490), .O(n500));
  nand2 g0437(.a(n412), .b(n410), .O(n501));
  nand2 g0438(.a(n412), .b(n407), .O(n502));
  nand2 g0439(.a(n410), .b(n407), .O(n503));
  and2  g0440(.a(n503), .b(n502), .O(n504));
  nand2 g0441(.a(n504), .b(n501), .O(n505));
  xor2  g0442(.a(n505), .b(n500), .O(n506));
  xor2  g0443(.a(n506), .b(n488), .O(n507));
  nand2 g0444(.a(n419), .b(n413), .O(n508));
  nand2 g0445(.a(n419), .b(n405), .O(n509));
  nand2 g0446(.a(n413), .b(n405), .O(n510));
  and2  g0447(.a(n510), .b(n509), .O(n511));
  nand2 g0448(.a(n511), .b(n508), .O(n512));
  xor2  g0449(.a(n512), .b(n507), .O(n513));
  xor2  g0450(.a(n513), .b(n486), .O(n514));
  nand2 g0451(.a(n426), .b(n420), .O(n515));
  nand2 g0452(.a(n426), .b(n403), .O(n516));
  nand2 g0453(.a(n420), .b(n403), .O(n517));
  and2  g0454(.a(n517), .b(n516), .O(n518));
  nand2 g0455(.a(n518), .b(n515), .O(n519));
  xor2  g0456(.a(n519), .b(n514), .O(n520));
  xor2  g0457(.a(n520), .b(n484), .O(n521));
  nand2 g0458(.a(n433), .b(n427), .O(n522));
  nand2 g0459(.a(n433), .b(n401), .O(n523));
  nand2 g0460(.a(n427), .b(n401), .O(n524));
  and2  g0461(.a(n524), .b(n523), .O(n525));
  nand2 g0462(.a(n525), .b(n522), .O(n526));
  xor2  g0463(.a(n526), .b(n521), .O(n527));
  xor2  g0464(.a(n527), .b(n482), .O(n528));
  nand2 g0465(.a(n440), .b(n434), .O(n529));
  nand2 g0466(.a(n440), .b(n399), .O(n530));
  nand2 g0467(.a(n434), .b(n399), .O(n531));
  and2  g0468(.a(n531), .b(n530), .O(n532));
  nand2 g0469(.a(n532), .b(n529), .O(n533));
  xor2  g0470(.a(n533), .b(n528), .O(n534));
  xor2  g0471(.a(n534), .b(n480), .O(n535));
  nand2 g0472(.a(n447), .b(n441), .O(n536));
  nand2 g0473(.a(n447), .b(n397), .O(n537));
  nand2 g0474(.a(n441), .b(n397), .O(n538));
  and2  g0475(.a(n538), .b(n537), .O(n539));
  nand2 g0476(.a(n539), .b(n536), .O(n540));
  xor2  g0477(.a(n540), .b(n535), .O(n541));
  xor2  g0478(.a(n541), .b(n478), .O(n542));
  nand2 g0479(.a(n455), .b(n448), .O(n543));
  nand2 g0480(.a(n455), .b(n395), .O(n544));
  nand2 g0481(.a(n448), .b(n395), .O(n545));
  and2  g0482(.a(n545), .b(n544), .O(n546));
  nand2 g0483(.a(n546), .b(n543), .O(n547));
  xor2  g0484(.a(n547), .b(n542), .O(n548));
  xor2  g0485(.a(n548), .b(n476), .O(n549));
  nand2 g0486(.a(n464), .b(n456), .O(n550));
  nand2 g0487(.a(n464), .b(n393), .O(n551));
  nand2 g0488(.a(n456), .b(n393), .O(n552));
  and2  g0489(.a(n552), .b(n551), .O(n553));
  nand2 g0490(.a(n553), .b(n550), .O(n554));
  xor2  g0491(.a(n554), .b(n549), .O(n555));
  xor2  g0492(.a(n555), .b(n474), .O(z11 ));
  nand2 g0493(.a(b12 ), .b(a0 ), .O(n557));
  inv1  g0494(.a(n557), .O(n558));
  nand2 g0495(.a(n555), .b(n473), .O(n559));
  nand2 g0496(.a(n473), .b(n468), .O(n560));
  nand2 g0497(.a(n555), .b(n468), .O(n561));
  and2  g0498(.a(n561), .b(n560), .O(n562));
  nand2 g0499(.a(n562), .b(n559), .O(n563));
  xor2  g0500(.a(n563), .b(n558), .O(n564));
  nand2 g0501(.a(b11 ), .b(a1 ), .O(n565));
  nand2 g0502(.a(b10 ), .b(a2 ), .O(n566));
  nand2 g0503(.a(b9 ), .b(a3 ), .O(n567));
  nand2 g0504(.a(b8 ), .b(a4 ), .O(n568));
  nand2 g0505(.a(b7 ), .b(a5 ), .O(n569));
  nand2 g0506(.a(b6 ), .b(a6 ), .O(n570));
  nand2 g0507(.a(b5 ), .b(a7 ), .O(n571));
  nand2 g0508(.a(b4 ), .b(a8 ), .O(n572));
  nand2 g0509(.a(b3 ), .b(a9 ), .O(n573));
  nand2 g0510(.a(b2 ), .b(a10 ), .O(n574));
  inv1  g0511(.a(n574), .O(n575));
  nand2 g0512(.a(b1 ), .b(a11 ), .O(n576));
  nand2 g0513(.a(b0 ), .b(a12 ), .O(n577));
  xor2  g0514(.a(n577), .b(n576), .O(n578));
  xor2  g0515(.a(n578), .b(n575), .O(n579));
  inv1  g0516(.a(n493), .O(n580));
  inv1  g0517(.a(n494), .O(n581));
  nand2 g0518(.a(n581), .b(n580), .O(n582));
  xor2  g0519(.a(n582), .b(n579), .O(n583));
  xor2  g0520(.a(n583), .b(n573), .O(n584));
  nand2 g0521(.a(n498), .b(n495), .O(n585));
  nand2 g0522(.a(n498), .b(n492), .O(n586));
  nand2 g0523(.a(n495), .b(n492), .O(n587));
  and2  g0524(.a(n587), .b(n586), .O(n588));
  nand2 g0525(.a(n588), .b(n585), .O(n589));
  xor2  g0526(.a(n589), .b(n584), .O(n590));
  xor2  g0527(.a(n590), .b(n572), .O(n591));
  nand2 g0528(.a(n505), .b(n499), .O(n592));
  nand2 g0529(.a(n505), .b(n490), .O(n593));
  nand2 g0530(.a(n499), .b(n490), .O(n594));
  and2  g0531(.a(n594), .b(n593), .O(n595));
  nand2 g0532(.a(n595), .b(n592), .O(n596));
  xor2  g0533(.a(n596), .b(n591), .O(n597));
  xor2  g0534(.a(n597), .b(n571), .O(n598));
  nand2 g0535(.a(n512), .b(n506), .O(n599));
  nand2 g0536(.a(n512), .b(n488), .O(n600));
  nand2 g0537(.a(n506), .b(n488), .O(n601));
  and2  g0538(.a(n601), .b(n600), .O(n602));
  nand2 g0539(.a(n602), .b(n599), .O(n603));
  xor2  g0540(.a(n603), .b(n598), .O(n604));
  xor2  g0541(.a(n604), .b(n570), .O(n605));
  nand2 g0542(.a(n519), .b(n513), .O(n606));
  nand2 g0543(.a(n519), .b(n486), .O(n607));
  nand2 g0544(.a(n513), .b(n486), .O(n608));
  and2  g0545(.a(n608), .b(n607), .O(n609));
  nand2 g0546(.a(n609), .b(n606), .O(n610));
  xor2  g0547(.a(n610), .b(n605), .O(n611));
  xor2  g0548(.a(n611), .b(n569), .O(n612));
  nand2 g0549(.a(n526), .b(n520), .O(n613));
  nand2 g0550(.a(n526), .b(n484), .O(n614));
  nand2 g0551(.a(n520), .b(n484), .O(n615));
  and2  g0552(.a(n615), .b(n614), .O(n616));
  nand2 g0553(.a(n616), .b(n613), .O(n617));
  xor2  g0554(.a(n617), .b(n612), .O(n618));
  xor2  g0555(.a(n618), .b(n568), .O(n619));
  nand2 g0556(.a(n533), .b(n527), .O(n620));
  nand2 g0557(.a(n533), .b(n482), .O(n621));
  nand2 g0558(.a(n527), .b(n482), .O(n622));
  and2  g0559(.a(n622), .b(n621), .O(n623));
  nand2 g0560(.a(n623), .b(n620), .O(n624));
  xor2  g0561(.a(n624), .b(n619), .O(n625));
  xor2  g0562(.a(n625), .b(n567), .O(n626));
  nand2 g0563(.a(n540), .b(n534), .O(n627));
  nand2 g0564(.a(n540), .b(n480), .O(n628));
  nand2 g0565(.a(n534), .b(n480), .O(n629));
  and2  g0566(.a(n629), .b(n628), .O(n630));
  nand2 g0567(.a(n630), .b(n627), .O(n631));
  xor2  g0568(.a(n631), .b(n626), .O(n632));
  xor2  g0569(.a(n632), .b(n566), .O(n633));
  nand2 g0570(.a(n547), .b(n541), .O(n634));
  nand2 g0571(.a(n547), .b(n478), .O(n635));
  nand2 g0572(.a(n541), .b(n478), .O(n636));
  and2  g0573(.a(n636), .b(n635), .O(n637));
  nand2 g0574(.a(n637), .b(n634), .O(n638));
  xor2  g0575(.a(n638), .b(n633), .O(n639));
  xor2  g0576(.a(n639), .b(n565), .O(n640));
  nand2 g0577(.a(n554), .b(n548), .O(n641));
  nand2 g0578(.a(n554), .b(n476), .O(n642));
  nand2 g0579(.a(n548), .b(n476), .O(n643));
  and2  g0580(.a(n643), .b(n642), .O(n644));
  nand2 g0581(.a(n644), .b(n641), .O(n645));
  xor2  g0582(.a(n645), .b(n640), .O(n646));
  xor2  g0583(.a(n646), .b(n564), .O(z12 ));
  nand2 g0584(.a(b13 ), .b(a0 ), .O(n648));
  inv1  g0585(.a(n648), .O(n649));
  nand2 g0586(.a(n646), .b(n563), .O(n650));
  nand2 g0587(.a(n563), .b(n558), .O(n651));
  nand2 g0588(.a(n646), .b(n558), .O(n652));
  and2  g0589(.a(n652), .b(n651), .O(n653));
  nand2 g0590(.a(n653), .b(n650), .O(n654));
  xor2  g0591(.a(n654), .b(n649), .O(n655));
  nand2 g0592(.a(b12 ), .b(a1 ), .O(n656));
  nand2 g0593(.a(b11 ), .b(a2 ), .O(n657));
  nand2 g0594(.a(b10 ), .b(a3 ), .O(n658));
  nand2 g0595(.a(b9 ), .b(a4 ), .O(n659));
  nand2 g0596(.a(b8 ), .b(a5 ), .O(n660));
  nand2 g0597(.a(b7 ), .b(a6 ), .O(n661));
  nand2 g0598(.a(b6 ), .b(a7 ), .O(n662));
  nand2 g0599(.a(b5 ), .b(a8 ), .O(n663));
  nand2 g0600(.a(b4 ), .b(a9 ), .O(n664));
  nand2 g0601(.a(b3 ), .b(a10 ), .O(n665));
  nand2 g0602(.a(b2 ), .b(a11 ), .O(n666));
  nand2 g0603(.a(b1 ), .b(a12 ), .O(n667));
  nand2 g0604(.a(b0 ), .b(a13 ), .O(n668));
  xor2  g0605(.a(n668), .b(n667), .O(n669));
  xor2  g0606(.a(n669), .b(n666), .O(n670));
  inv1  g0607(.a(n576), .O(n671));
  inv1  g0608(.a(n577), .O(n672));
  nand2 g0609(.a(n672), .b(n671), .O(n673));
  xor2  g0610(.a(n673), .b(n670), .O(n674));
  xor2  g0611(.a(n674), .b(n665), .O(n675));
  inv1  g0612(.a(n582), .O(n676));
  nand2 g0613(.a(n676), .b(n578), .O(n677));
  nand2 g0614(.a(n676), .b(n575), .O(n678));
  nand2 g0615(.a(n578), .b(n575), .O(n679));
  and2  g0616(.a(n679), .b(n678), .O(n680));
  nand2 g0617(.a(n680), .b(n677), .O(n681));
  xor2  g0618(.a(n681), .b(n675), .O(n682));
  xor2  g0619(.a(n682), .b(n664), .O(n683));
  inv1  g0620(.a(n583), .O(n684));
  nand2 g0621(.a(n589), .b(n684), .O(n685));
  inv1  g0622(.a(n573), .O(n686));
  nand2 g0623(.a(n589), .b(n686), .O(n687));
  nand2 g0624(.a(n684), .b(n686), .O(n688));
  and2  g0625(.a(n688), .b(n687), .O(n689));
  nand2 g0626(.a(n689), .b(n685), .O(n690));
  xor2  g0627(.a(n690), .b(n683), .O(n691));
  xor2  g0628(.a(n691), .b(n663), .O(n692));
  nand2 g0629(.a(n596), .b(n590), .O(n693));
  inv1  g0630(.a(n572), .O(n694));
  nand2 g0631(.a(n596), .b(n694), .O(n695));
  nand2 g0632(.a(n590), .b(n694), .O(n696));
  and2  g0633(.a(n696), .b(n695), .O(n697));
  nand2 g0634(.a(n697), .b(n693), .O(n698));
  xor2  g0635(.a(n698), .b(n692), .O(n699));
  xor2  g0636(.a(n699), .b(n662), .O(n700));
  inv1  g0637(.a(n597), .O(n701));
  nand2 g0638(.a(n603), .b(n701), .O(n702));
  inv1  g0639(.a(n571), .O(n703));
  nand2 g0640(.a(n603), .b(n703), .O(n704));
  nand2 g0641(.a(n701), .b(n703), .O(n705));
  and2  g0642(.a(n705), .b(n704), .O(n706));
  nand2 g0643(.a(n706), .b(n702), .O(n707));
  xor2  g0644(.a(n707), .b(n700), .O(n708));
  xor2  g0645(.a(n708), .b(n661), .O(n709));
  nand2 g0646(.a(n610), .b(n604), .O(n710));
  inv1  g0647(.a(n570), .O(n711));
  nand2 g0648(.a(n610), .b(n711), .O(n712));
  nand2 g0649(.a(n604), .b(n711), .O(n713));
  and2  g0650(.a(n713), .b(n712), .O(n714));
  nand2 g0651(.a(n714), .b(n710), .O(n715));
  xor2  g0652(.a(n715), .b(n709), .O(n716));
  xor2  g0653(.a(n716), .b(n660), .O(n717));
  inv1  g0654(.a(n611), .O(n718));
  nand2 g0655(.a(n617), .b(n718), .O(n719));
  inv1  g0656(.a(n569), .O(n720));
  nand2 g0657(.a(n617), .b(n720), .O(n721));
  nand2 g0658(.a(n718), .b(n720), .O(n722));
  and2  g0659(.a(n722), .b(n721), .O(n723));
  nand2 g0660(.a(n723), .b(n719), .O(n724));
  xor2  g0661(.a(n724), .b(n717), .O(n725));
  xor2  g0662(.a(n725), .b(n659), .O(n726));
  nand2 g0663(.a(n624), .b(n618), .O(n727));
  inv1  g0664(.a(n568), .O(n728));
  nand2 g0665(.a(n624), .b(n728), .O(n729));
  nand2 g0666(.a(n618), .b(n728), .O(n730));
  and2  g0667(.a(n730), .b(n729), .O(n731));
  nand2 g0668(.a(n731), .b(n727), .O(n732));
  xor2  g0669(.a(n732), .b(n726), .O(n733));
  xor2  g0670(.a(n733), .b(n658), .O(n734));
  inv1  g0671(.a(n625), .O(n735));
  nand2 g0672(.a(n631), .b(n735), .O(n736));
  inv1  g0673(.a(n567), .O(n737));
  nand2 g0674(.a(n631), .b(n737), .O(n738));
  nand2 g0675(.a(n735), .b(n737), .O(n739));
  and2  g0676(.a(n739), .b(n738), .O(n740));
  nand2 g0677(.a(n740), .b(n736), .O(n741));
  xor2  g0678(.a(n741), .b(n734), .O(n742));
  xor2  g0679(.a(n742), .b(n657), .O(n743));
  nand2 g0680(.a(n638), .b(n632), .O(n744));
  inv1  g0681(.a(n566), .O(n745));
  nand2 g0682(.a(n638), .b(n745), .O(n746));
  nand2 g0683(.a(n632), .b(n745), .O(n747));
  and2  g0684(.a(n747), .b(n746), .O(n748));
  nand2 g0685(.a(n748), .b(n744), .O(n749));
  xor2  g0686(.a(n749), .b(n743), .O(n750));
  xor2  g0687(.a(n750), .b(n656), .O(n751));
  inv1  g0688(.a(n639), .O(n752));
  nand2 g0689(.a(n645), .b(n752), .O(n753));
  inv1  g0690(.a(n565), .O(n754));
  nand2 g0691(.a(n645), .b(n754), .O(n755));
  nand2 g0692(.a(n752), .b(n754), .O(n756));
  and2  g0693(.a(n756), .b(n755), .O(n757));
  nand2 g0694(.a(n757), .b(n753), .O(n758));
  xor2  g0695(.a(n758), .b(n751), .O(n759));
  xor2  g0696(.a(n759), .b(n655), .O(z13 ));
  nand2 g0697(.a(b14 ), .b(a0 ), .O(n761));
  inv1  g0698(.a(n761), .O(n762));
  nand2 g0699(.a(n759), .b(n654), .O(n763));
  nand2 g0700(.a(n654), .b(n649), .O(n764));
  nand2 g0701(.a(n759), .b(n649), .O(n765));
  and2  g0702(.a(n765), .b(n764), .O(n766));
  nand2 g0703(.a(n766), .b(n763), .O(n767));
  xor2  g0704(.a(n767), .b(n762), .O(n768));
  nand2 g0705(.a(b13 ), .b(a1 ), .O(n769));
  nand2 g0706(.a(b12 ), .b(a2 ), .O(n770));
  nand2 g0707(.a(b11 ), .b(a3 ), .O(n771));
  nand2 g0708(.a(b10 ), .b(a4 ), .O(n772));
  nand2 g0709(.a(b9 ), .b(a5 ), .O(n773));
  nand2 g0710(.a(b8 ), .b(a6 ), .O(n774));
  nand2 g0711(.a(b7 ), .b(a7 ), .O(n775));
  nand2 g0712(.a(b6 ), .b(a8 ), .O(n776));
  nand2 g0713(.a(b5 ), .b(a9 ), .O(n777));
  nand2 g0714(.a(b4 ), .b(a10 ), .O(n778));
  nand2 g0715(.a(b3 ), .b(a11 ), .O(n779));
  nand2 g0716(.a(b2 ), .b(a12 ), .O(n780));
  inv1  g0717(.a(n780), .O(n781));
  nand2 g0718(.a(b1 ), .b(a13 ), .O(n782));
  nand2 g0719(.a(b0 ), .b(a14 ), .O(n783));
  xor2  g0720(.a(n783), .b(n782), .O(n784));
  xor2  g0721(.a(n784), .b(n781), .O(n785));
  inv1  g0722(.a(n667), .O(n786));
  inv1  g0723(.a(n668), .O(n787));
  nand2 g0724(.a(n787), .b(n786), .O(n788));
  xor2  g0725(.a(n788), .b(n785), .O(n789));
  xor2  g0726(.a(n789), .b(n779), .O(n790));
  inv1  g0727(.a(n673), .O(n791));
  nand2 g0728(.a(n791), .b(n669), .O(n792));
  inv1  g0729(.a(n666), .O(n793));
  nand2 g0730(.a(n791), .b(n793), .O(n794));
  nand2 g0731(.a(n669), .b(n793), .O(n795));
  and2  g0732(.a(n795), .b(n794), .O(n796));
  nand2 g0733(.a(n796), .b(n792), .O(n797));
  xor2  g0734(.a(n797), .b(n790), .O(n798));
  xor2  g0735(.a(n798), .b(n778), .O(n799));
  nand2 g0736(.a(n681), .b(n674), .O(n800));
  inv1  g0737(.a(n665), .O(n801));
  nand2 g0738(.a(n681), .b(n801), .O(n802));
  nand2 g0739(.a(n674), .b(n801), .O(n803));
  and2  g0740(.a(n803), .b(n802), .O(n804));
  nand2 g0741(.a(n804), .b(n800), .O(n805));
  xor2  g0742(.a(n805), .b(n799), .O(n806));
  xor2  g0743(.a(n806), .b(n777), .O(n807));
  inv1  g0744(.a(n682), .O(n808));
  nand2 g0745(.a(n690), .b(n808), .O(n809));
  inv1  g0746(.a(n664), .O(n810));
  nand2 g0747(.a(n690), .b(n810), .O(n811));
  nand2 g0748(.a(n808), .b(n810), .O(n812));
  and2  g0749(.a(n812), .b(n811), .O(n813));
  nand2 g0750(.a(n813), .b(n809), .O(n814));
  xor2  g0751(.a(n814), .b(n807), .O(n815));
  xor2  g0752(.a(n815), .b(n776), .O(n816));
  nand2 g0753(.a(n698), .b(n691), .O(n817));
  inv1  g0754(.a(n663), .O(n818));
  nand2 g0755(.a(n698), .b(n818), .O(n819));
  nand2 g0756(.a(n691), .b(n818), .O(n820));
  and2  g0757(.a(n820), .b(n819), .O(n821));
  nand2 g0758(.a(n821), .b(n817), .O(n822));
  xor2  g0759(.a(n822), .b(n816), .O(n823));
  xor2  g0760(.a(n823), .b(n775), .O(n824));
  inv1  g0761(.a(n699), .O(n825));
  nand2 g0762(.a(n707), .b(n825), .O(n826));
  inv1  g0763(.a(n662), .O(n827));
  nand2 g0764(.a(n707), .b(n827), .O(n828));
  nand2 g0765(.a(n825), .b(n827), .O(n829));
  and2  g0766(.a(n829), .b(n828), .O(n830));
  nand2 g0767(.a(n830), .b(n826), .O(n831));
  xor2  g0768(.a(n831), .b(n824), .O(n832));
  xor2  g0769(.a(n832), .b(n774), .O(n833));
  nand2 g0770(.a(n715), .b(n708), .O(n834));
  inv1  g0771(.a(n661), .O(n835));
  nand2 g0772(.a(n715), .b(n835), .O(n836));
  nand2 g0773(.a(n708), .b(n835), .O(n837));
  and2  g0774(.a(n837), .b(n836), .O(n838));
  nand2 g0775(.a(n838), .b(n834), .O(n839));
  xor2  g0776(.a(n839), .b(n833), .O(n840));
  xor2  g0777(.a(n840), .b(n773), .O(n841));
  inv1  g0778(.a(n716), .O(n842));
  nand2 g0779(.a(n724), .b(n842), .O(n843));
  inv1  g0780(.a(n660), .O(n844));
  nand2 g0781(.a(n724), .b(n844), .O(n845));
  nand2 g0782(.a(n842), .b(n844), .O(n846));
  and2  g0783(.a(n846), .b(n845), .O(n847));
  nand2 g0784(.a(n847), .b(n843), .O(n848));
  xor2  g0785(.a(n848), .b(n841), .O(n849));
  xor2  g0786(.a(n849), .b(n772), .O(n850));
  nand2 g0787(.a(n732), .b(n725), .O(n851));
  inv1  g0788(.a(n659), .O(n852));
  nand2 g0789(.a(n732), .b(n852), .O(n853));
  nand2 g0790(.a(n725), .b(n852), .O(n854));
  and2  g0791(.a(n854), .b(n853), .O(n855));
  nand2 g0792(.a(n855), .b(n851), .O(n856));
  xor2  g0793(.a(n856), .b(n850), .O(n857));
  xor2  g0794(.a(n857), .b(n771), .O(n858));
  inv1  g0795(.a(n733), .O(n859));
  nand2 g0796(.a(n741), .b(n859), .O(n860));
  inv1  g0797(.a(n658), .O(n861));
  nand2 g0798(.a(n741), .b(n861), .O(n862));
  nand2 g0799(.a(n859), .b(n861), .O(n863));
  and2  g0800(.a(n863), .b(n862), .O(n864));
  nand2 g0801(.a(n864), .b(n860), .O(n865));
  xor2  g0802(.a(n865), .b(n858), .O(n866));
  xor2  g0803(.a(n866), .b(n770), .O(n867));
  nand2 g0804(.a(n749), .b(n742), .O(n868));
  inv1  g0805(.a(n657), .O(n869));
  nand2 g0806(.a(n749), .b(n869), .O(n870));
  nand2 g0807(.a(n742), .b(n869), .O(n871));
  and2  g0808(.a(n871), .b(n870), .O(n872));
  nand2 g0809(.a(n872), .b(n868), .O(n873));
  xor2  g0810(.a(n873), .b(n867), .O(n874));
  xor2  g0811(.a(n874), .b(n769), .O(n875));
  inv1  g0812(.a(n750), .O(n876));
  nand2 g0813(.a(n758), .b(n876), .O(n877));
  inv1  g0814(.a(n656), .O(n878));
  nand2 g0815(.a(n758), .b(n878), .O(n879));
  nand2 g0816(.a(n876), .b(n878), .O(n880));
  and2  g0817(.a(n880), .b(n879), .O(n881));
  nand2 g0818(.a(n881), .b(n877), .O(n882));
  xor2  g0819(.a(n882), .b(n875), .O(n883));
  xor2  g0820(.a(n883), .b(n768), .O(z14 ));
  nand2 g0821(.a(b15 ), .b(a0 ), .O(n885));
  inv1  g0822(.a(n885), .O(n886));
  nand2 g0823(.a(n883), .b(n767), .O(n887));
  nand2 g0824(.a(n767), .b(n762), .O(n888));
  nand2 g0825(.a(n883), .b(n762), .O(n889));
  and2  g0826(.a(n889), .b(n888), .O(n890));
  nand2 g0827(.a(n890), .b(n887), .O(n891));
  xor2  g0828(.a(n891), .b(n886), .O(n892));
  nand2 g0829(.a(b14 ), .b(a1 ), .O(n893));
  nand2 g0830(.a(b13 ), .b(a2 ), .O(n894));
  nand2 g0831(.a(b12 ), .b(a3 ), .O(n895));
  nand2 g0832(.a(b11 ), .b(a4 ), .O(n896));
  nand2 g0833(.a(b10 ), .b(a5 ), .O(n897));
  nand2 g0834(.a(b9 ), .b(a6 ), .O(n898));
  nand2 g0835(.a(b8 ), .b(a7 ), .O(n899));
  nand2 g0836(.a(b7 ), .b(a8 ), .O(n900));
  nand2 g0837(.a(b6 ), .b(a9 ), .O(n901));
  nand2 g0838(.a(b5 ), .b(a10 ), .O(n902));
  nand2 g0839(.a(b4 ), .b(a11 ), .O(n903));
  nand2 g0840(.a(b3 ), .b(a12 ), .O(n904));
  nand2 g0841(.a(b2 ), .b(a13 ), .O(n905));
  nand2 g0842(.a(b1 ), .b(a14 ), .O(n906));
  nand2 g0843(.a(b0 ), .b(a15 ), .O(n907));
  xor2  g0844(.a(n907), .b(n906), .O(n908));
  xor2  g0845(.a(n908), .b(n905), .O(n909));
  inv1  g0846(.a(n782), .O(n910));
  inv1  g0847(.a(n783), .O(n911));
  nand2 g0848(.a(n911), .b(n910), .O(n912));
  xor2  g0849(.a(n912), .b(n909), .O(n913));
  xor2  g0850(.a(n913), .b(n904), .O(n914));
  inv1  g0851(.a(n788), .O(n915));
  nand2 g0852(.a(n915), .b(n784), .O(n916));
  nand2 g0853(.a(n915), .b(n781), .O(n917));
  nand2 g0854(.a(n784), .b(n781), .O(n918));
  and2  g0855(.a(n918), .b(n917), .O(n919));
  nand2 g0856(.a(n919), .b(n916), .O(n920));
  xor2  g0857(.a(n920), .b(n914), .O(n921));
  xor2  g0858(.a(n921), .b(n903), .O(n922));
  inv1  g0859(.a(n789), .O(n923));
  nand2 g0860(.a(n797), .b(n923), .O(n924));
  inv1  g0861(.a(n779), .O(n925));
  nand2 g0862(.a(n797), .b(n925), .O(n926));
  nand2 g0863(.a(n923), .b(n925), .O(n927));
  and2  g0864(.a(n927), .b(n926), .O(n928));
  nand2 g0865(.a(n928), .b(n924), .O(n929));
  xor2  g0866(.a(n929), .b(n922), .O(n930));
  xor2  g0867(.a(n930), .b(n902), .O(n931));
  nand2 g0868(.a(n805), .b(n798), .O(n932));
  inv1  g0869(.a(n778), .O(n933));
  nand2 g0870(.a(n805), .b(n933), .O(n934));
  nand2 g0871(.a(n798), .b(n933), .O(n935));
  and2  g0872(.a(n935), .b(n934), .O(n936));
  nand2 g0873(.a(n936), .b(n932), .O(n937));
  xor2  g0874(.a(n937), .b(n931), .O(n938));
  xor2  g0875(.a(n938), .b(n901), .O(n939));
  inv1  g0876(.a(n806), .O(n940));
  nand2 g0877(.a(n814), .b(n940), .O(n941));
  inv1  g0878(.a(n777), .O(n942));
  nand2 g0879(.a(n814), .b(n942), .O(n943));
  nand2 g0880(.a(n940), .b(n942), .O(n944));
  and2  g0881(.a(n944), .b(n943), .O(n945));
  nand2 g0882(.a(n945), .b(n941), .O(n946));
  xor2  g0883(.a(n946), .b(n939), .O(n947));
  xor2  g0884(.a(n947), .b(n900), .O(n948));
  nand2 g0885(.a(n822), .b(n815), .O(n949));
  inv1  g0886(.a(n776), .O(n950));
  nand2 g0887(.a(n822), .b(n950), .O(n951));
  nand2 g0888(.a(n815), .b(n950), .O(n952));
  and2  g0889(.a(n952), .b(n951), .O(n953));
  nand2 g0890(.a(n953), .b(n949), .O(n954));
  xor2  g0891(.a(n954), .b(n948), .O(n955));
  xor2  g0892(.a(n955), .b(n899), .O(n956));
  inv1  g0893(.a(n823), .O(n957));
  nand2 g0894(.a(n831), .b(n957), .O(n958));
  inv1  g0895(.a(n775), .O(n959));
  nand2 g0896(.a(n831), .b(n959), .O(n960));
  nand2 g0897(.a(n957), .b(n959), .O(n961));
  and2  g0898(.a(n961), .b(n960), .O(n962));
  nand2 g0899(.a(n962), .b(n958), .O(n963));
  xor2  g0900(.a(n963), .b(n956), .O(n964));
  xor2  g0901(.a(n964), .b(n898), .O(n965));
  nand2 g0902(.a(n839), .b(n832), .O(n966));
  inv1  g0903(.a(n774), .O(n967));
  nand2 g0904(.a(n839), .b(n967), .O(n968));
  nand2 g0905(.a(n832), .b(n967), .O(n969));
  and2  g0906(.a(n969), .b(n968), .O(n970));
  nand2 g0907(.a(n970), .b(n966), .O(n971));
  xor2  g0908(.a(n971), .b(n965), .O(n972));
  xor2  g0909(.a(n972), .b(n897), .O(n973));
  inv1  g0910(.a(n840), .O(n974));
  nand2 g0911(.a(n848), .b(n974), .O(n975));
  inv1  g0912(.a(n773), .O(n976));
  nand2 g0913(.a(n848), .b(n976), .O(n977));
  nand2 g0914(.a(n974), .b(n976), .O(n978));
  and2  g0915(.a(n978), .b(n977), .O(n979));
  nand2 g0916(.a(n979), .b(n975), .O(n980));
  xor2  g0917(.a(n980), .b(n973), .O(n981));
  xor2  g0918(.a(n981), .b(n896), .O(n982));
  nand2 g0919(.a(n856), .b(n849), .O(n983));
  inv1  g0920(.a(n772), .O(n984));
  nand2 g0921(.a(n856), .b(n984), .O(n985));
  nand2 g0922(.a(n849), .b(n984), .O(n986));
  and2  g0923(.a(n986), .b(n985), .O(n987));
  nand2 g0924(.a(n987), .b(n983), .O(n988));
  xor2  g0925(.a(n988), .b(n982), .O(n989));
  xor2  g0926(.a(n989), .b(n895), .O(n990));
  inv1  g0927(.a(n857), .O(n991));
  nand2 g0928(.a(n865), .b(n991), .O(n992));
  inv1  g0929(.a(n771), .O(n993));
  nand2 g0930(.a(n865), .b(n993), .O(n994));
  nand2 g0931(.a(n991), .b(n993), .O(n995));
  and2  g0932(.a(n995), .b(n994), .O(n996));
  nand2 g0933(.a(n996), .b(n992), .O(n997));
  xor2  g0934(.a(n997), .b(n990), .O(n998));
  xor2  g0935(.a(n998), .b(n894), .O(n999));
  nand2 g0936(.a(n873), .b(n866), .O(n1000));
  inv1  g0937(.a(n770), .O(n1001));
  nand2 g0938(.a(n873), .b(n1001), .O(n1002));
  nand2 g0939(.a(n866), .b(n1001), .O(n1003));
  and2  g0940(.a(n1003), .b(n1002), .O(n1004));
  nand2 g0941(.a(n1004), .b(n1000), .O(n1005));
  xor2  g0942(.a(n1005), .b(n999), .O(n1006));
  xor2  g0943(.a(n1006), .b(n893), .O(n1007));
  inv1  g0944(.a(n874), .O(n1008));
  nand2 g0945(.a(n882), .b(n1008), .O(n1009));
  inv1  g0946(.a(n769), .O(n1010));
  nand2 g0947(.a(n882), .b(n1010), .O(n1011));
  nand2 g0948(.a(n1008), .b(n1010), .O(n1012));
  and2  g0949(.a(n1012), .b(n1011), .O(n1013));
  nand2 g0950(.a(n1013), .b(n1009), .O(n1014));
  xor2  g0951(.a(n1014), .b(n1007), .O(n1015));
  xor2  g0952(.a(n1015), .b(n892), .O(z15 ));
  nand2 g0953(.a(b15 ), .b(a1 ), .O(n1017));
  nand2 g0954(.a(b14 ), .b(a2 ), .O(n1018));
  nand2 g0955(.a(b13 ), .b(a3 ), .O(n1019));
  nand2 g0956(.a(b12 ), .b(a4 ), .O(n1020));
  nand2 g0957(.a(b11 ), .b(a5 ), .O(n1021));
  nand2 g0958(.a(b10 ), .b(a6 ), .O(n1022));
  nand2 g0959(.a(b9 ), .b(a7 ), .O(n1023));
  nand2 g0960(.a(b8 ), .b(a8 ), .O(n1024));
  nand2 g0961(.a(b7 ), .b(a9 ), .O(n1025));
  nand2 g0962(.a(b6 ), .b(a10 ), .O(n1026));
  nand2 g0963(.a(b5 ), .b(a11 ), .O(n1027));
  nand2 g0964(.a(b4 ), .b(a12 ), .O(n1028));
  nand2 g0965(.a(b3 ), .b(a13 ), .O(n1029));
  inv1  g0966(.a(n1029), .O(n1030));
  nand2 g0967(.a(b2 ), .b(a14 ), .O(n1031));
  nand2 g0968(.a(b1 ), .b(a15 ), .O(n1032));
  xnor2 g0969(.a(n1032), .b(n1031), .O(n1033));
  inv1  g0970(.a(n906), .O(n1034));
  inv1  g0971(.a(n907), .O(n1035));
  nand2 g0972(.a(n1035), .b(n1034), .O(n1036));
  xnor2 g0973(.a(n1036), .b(n1033), .O(n1037));
  xor2  g0974(.a(n1037), .b(n1030), .O(n1038));
  inv1  g0975(.a(n912), .O(n1039));
  nand2 g0976(.a(n1039), .b(n908), .O(n1040));
  inv1  g0977(.a(n905), .O(n1041));
  nand2 g0978(.a(n1039), .b(n1041), .O(n1042));
  nand2 g0979(.a(n908), .b(n1041), .O(n1043));
  and2  g0980(.a(n1043), .b(n1042), .O(n1044));
  nand2 g0981(.a(n1044), .b(n1040), .O(n1045));
  xnor2 g0982(.a(n1045), .b(n1038), .O(n1046));
  xor2  g0983(.a(n1046), .b(n1028), .O(n1047));
  nand2 g0984(.a(n920), .b(n913), .O(n1048));
  inv1  g0985(.a(n904), .O(n1049));
  nand2 g0986(.a(n920), .b(n1049), .O(n1050));
  nand2 g0987(.a(n913), .b(n1049), .O(n1051));
  and2  g0988(.a(n1051), .b(n1050), .O(n1052));
  nand2 g0989(.a(n1052), .b(n1048), .O(n1053));
  xor2  g0990(.a(n1053), .b(n1047), .O(n1054));
  xor2  g0991(.a(n1054), .b(n1027), .O(n1055));
  inv1  g0992(.a(n921), .O(n1056));
  nand2 g0993(.a(n929), .b(n1056), .O(n1057));
  inv1  g0994(.a(n903), .O(n1058));
  nand2 g0995(.a(n929), .b(n1058), .O(n1059));
  nand2 g0996(.a(n1056), .b(n1058), .O(n1060));
  and2  g0997(.a(n1060), .b(n1059), .O(n1061));
  nand2 g0998(.a(n1061), .b(n1057), .O(n1062));
  xor2  g0999(.a(n1062), .b(n1055), .O(n1063));
  xor2  g1000(.a(n1063), .b(n1026), .O(n1064));
  nand2 g1001(.a(n937), .b(n930), .O(n1065));
  inv1  g1002(.a(n902), .O(n1066));
  nand2 g1003(.a(n937), .b(n1066), .O(n1067));
  nand2 g1004(.a(n930), .b(n1066), .O(n1068));
  and2  g1005(.a(n1068), .b(n1067), .O(n1069));
  nand2 g1006(.a(n1069), .b(n1065), .O(n1070));
  xor2  g1007(.a(n1070), .b(n1064), .O(n1071));
  xor2  g1008(.a(n1071), .b(n1025), .O(n1072));
  inv1  g1009(.a(n938), .O(n1073));
  nand2 g1010(.a(n946), .b(n1073), .O(n1074));
  inv1  g1011(.a(n901), .O(n1075));
  nand2 g1012(.a(n946), .b(n1075), .O(n1076));
  nand2 g1013(.a(n1073), .b(n1075), .O(n1077));
  and2  g1014(.a(n1077), .b(n1076), .O(n1078));
  nand2 g1015(.a(n1078), .b(n1074), .O(n1079));
  xor2  g1016(.a(n1079), .b(n1072), .O(n1080));
  xor2  g1017(.a(n1080), .b(n1024), .O(n1081));
  nand2 g1018(.a(n954), .b(n947), .O(n1082));
  inv1  g1019(.a(n900), .O(n1083));
  nand2 g1020(.a(n954), .b(n1083), .O(n1084));
  nand2 g1021(.a(n947), .b(n1083), .O(n1085));
  and2  g1022(.a(n1085), .b(n1084), .O(n1086));
  nand2 g1023(.a(n1086), .b(n1082), .O(n1087));
  xor2  g1024(.a(n1087), .b(n1081), .O(n1088));
  xor2  g1025(.a(n1088), .b(n1023), .O(n1089));
  inv1  g1026(.a(n955), .O(n1090));
  nand2 g1027(.a(n963), .b(n1090), .O(n1091));
  inv1  g1028(.a(n899), .O(n1092));
  nand2 g1029(.a(n963), .b(n1092), .O(n1093));
  nand2 g1030(.a(n1090), .b(n1092), .O(n1094));
  and2  g1031(.a(n1094), .b(n1093), .O(n1095));
  nand2 g1032(.a(n1095), .b(n1091), .O(n1096));
  xor2  g1033(.a(n1096), .b(n1089), .O(n1097));
  xor2  g1034(.a(n1097), .b(n1022), .O(n1098));
  nand2 g1035(.a(n971), .b(n964), .O(n1099));
  inv1  g1036(.a(n898), .O(n1100));
  nand2 g1037(.a(n971), .b(n1100), .O(n1101));
  nand2 g1038(.a(n964), .b(n1100), .O(n1102));
  and2  g1039(.a(n1102), .b(n1101), .O(n1103));
  nand2 g1040(.a(n1103), .b(n1099), .O(n1104));
  xor2  g1041(.a(n1104), .b(n1098), .O(n1105));
  xor2  g1042(.a(n1105), .b(n1021), .O(n1106));
  inv1  g1043(.a(n972), .O(n1107));
  nand2 g1044(.a(n980), .b(n1107), .O(n1108));
  inv1  g1045(.a(n897), .O(n1109));
  nand2 g1046(.a(n980), .b(n1109), .O(n1110));
  nand2 g1047(.a(n1107), .b(n1109), .O(n1111));
  and2  g1048(.a(n1111), .b(n1110), .O(n1112));
  nand2 g1049(.a(n1112), .b(n1108), .O(n1113));
  xor2  g1050(.a(n1113), .b(n1106), .O(n1114));
  xor2  g1051(.a(n1114), .b(n1020), .O(n1115));
  nand2 g1052(.a(n988), .b(n981), .O(n1116));
  inv1  g1053(.a(n896), .O(n1117));
  nand2 g1054(.a(n988), .b(n1117), .O(n1118));
  nand2 g1055(.a(n981), .b(n1117), .O(n1119));
  and2  g1056(.a(n1119), .b(n1118), .O(n1120));
  nand2 g1057(.a(n1120), .b(n1116), .O(n1121));
  xor2  g1058(.a(n1121), .b(n1115), .O(n1122));
  xor2  g1059(.a(n1122), .b(n1019), .O(n1123));
  inv1  g1060(.a(n989), .O(n1124));
  nand2 g1061(.a(n997), .b(n1124), .O(n1125));
  inv1  g1062(.a(n895), .O(n1126));
  nand2 g1063(.a(n997), .b(n1126), .O(n1127));
  nand2 g1064(.a(n1124), .b(n1126), .O(n1128));
  and2  g1065(.a(n1128), .b(n1127), .O(n1129));
  nand2 g1066(.a(n1129), .b(n1125), .O(n1130));
  xor2  g1067(.a(n1130), .b(n1123), .O(n1131));
  xor2  g1068(.a(n1131), .b(n1018), .O(n1132));
  nand2 g1069(.a(n1005), .b(n998), .O(n1133));
  inv1  g1070(.a(n894), .O(n1134));
  nand2 g1071(.a(n1005), .b(n1134), .O(n1135));
  nand2 g1072(.a(n998), .b(n1134), .O(n1136));
  and2  g1073(.a(n1136), .b(n1135), .O(n1137));
  nand2 g1074(.a(n1137), .b(n1133), .O(n1138));
  xor2  g1075(.a(n1138), .b(n1132), .O(n1139));
  xor2  g1076(.a(n1139), .b(n1017), .O(n1140));
  inv1  g1077(.a(n1006), .O(n1141));
  nand2 g1078(.a(n1014), .b(n1141), .O(n1142));
  inv1  g1079(.a(n893), .O(n1143));
  nand2 g1080(.a(n1014), .b(n1143), .O(n1144));
  nand2 g1081(.a(n1141), .b(n1143), .O(n1145));
  and2  g1082(.a(n1145), .b(n1144), .O(n1146));
  nand2 g1083(.a(n1146), .b(n1142), .O(n1147));
  xor2  g1084(.a(n1147), .b(n1140), .O(n1148));
  nand2 g1085(.a(n1015), .b(n891), .O(n1149));
  nand2 g1086(.a(n891), .b(n886), .O(n1150));
  nand2 g1087(.a(n1015), .b(n886), .O(n1151));
  and2  g1088(.a(n1151), .b(n1150), .O(n1152));
  nand2 g1089(.a(n1152), .b(n1149), .O(n1153));
  xor2  g1090(.a(n1153), .b(n1148), .O(z16 ));
  and2  g1091(.a(n1153), .b(n1148), .O(n1155));
  nand2 g1092(.a(b15 ), .b(a2 ), .O(n1156));
  inv1  g1093(.a(n1156), .O(n1157));
  nand2 g1094(.a(b14 ), .b(a3 ), .O(n1158));
  inv1  g1095(.a(n1158), .O(n1159));
  nand2 g1096(.a(b13 ), .b(a4 ), .O(n1160));
  inv1  g1097(.a(n1160), .O(n1161));
  nand2 g1098(.a(b12 ), .b(a5 ), .O(n1162));
  inv1  g1099(.a(n1162), .O(n1163));
  nand2 g1100(.a(b11 ), .b(a6 ), .O(n1164));
  inv1  g1101(.a(n1164), .O(n1165));
  nand2 g1102(.a(b10 ), .b(a7 ), .O(n1166));
  inv1  g1103(.a(n1166), .O(n1167));
  nand2 g1104(.a(b9 ), .b(a8 ), .O(n1168));
  inv1  g1105(.a(n1168), .O(n1169));
  nand2 g1106(.a(b8 ), .b(a9 ), .O(n1170));
  inv1  g1107(.a(n1170), .O(n1171));
  nand2 g1108(.a(b7 ), .b(a10 ), .O(n1172));
  inv1  g1109(.a(n1172), .O(n1173));
  nand2 g1110(.a(b6 ), .b(a11 ), .O(n1174));
  inv1  g1111(.a(n1174), .O(n1175));
  nand2 g1112(.a(b5 ), .b(a12 ), .O(n1176));
  inv1  g1113(.a(n1176), .O(n1177));
  nand2 g1114(.a(b4 ), .b(a13 ), .O(n1178));
  inv1  g1115(.a(n1178), .O(n1179));
  nand2 g1116(.a(b3 ), .b(a14 ), .O(n1180));
  nand2 g1117(.a(b2 ), .b(a15 ), .O(n1181));
  xnor2 g1118(.a(n1181), .b(n1180), .O(n1182));
  inv1  g1119(.a(n1032), .O(n1183));
  inv1  g1120(.a(n1036), .O(n1184));
  nand2 g1121(.a(n1184), .b(n1183), .O(n1185));
  inv1  g1122(.a(n1031), .O(n1186));
  nand2 g1123(.a(n1184), .b(n1186), .O(n1187));
  nand2 g1124(.a(n1183), .b(n1186), .O(n1188));
  and2  g1125(.a(n1188), .b(n1187), .O(n1189));
  nand2 g1126(.a(n1189), .b(n1185), .O(n1190));
  xor2  g1127(.a(n1190), .b(n1182), .O(n1191));
  xor2  g1128(.a(n1191), .b(n1179), .O(n1192));
  inv1  g1129(.a(n1037), .O(n1193));
  nand2 g1130(.a(n1045), .b(n1193), .O(n1194));
  nand2 g1131(.a(n1045), .b(n1030), .O(n1195));
  nand2 g1132(.a(n1193), .b(n1030), .O(n1196));
  and2  g1133(.a(n1196), .b(n1195), .O(n1197));
  nand2 g1134(.a(n1197), .b(n1194), .O(n1198));
  xor2  g1135(.a(n1198), .b(n1192), .O(n1199));
  xor2  g1136(.a(n1199), .b(n1177), .O(n1200));
  nand2 g1137(.a(n1053), .b(n1046), .O(n1201));
  inv1  g1138(.a(n1028), .O(n1202));
  nand2 g1139(.a(n1053), .b(n1202), .O(n1203));
  nand2 g1140(.a(n1046), .b(n1202), .O(n1204));
  and2  g1141(.a(n1204), .b(n1203), .O(n1205));
  nand2 g1142(.a(n1205), .b(n1201), .O(n1206));
  xor2  g1143(.a(n1206), .b(n1200), .O(n1207));
  xor2  g1144(.a(n1207), .b(n1175), .O(n1208));
  inv1  g1145(.a(n1054), .O(n1209));
  nand2 g1146(.a(n1062), .b(n1209), .O(n1210));
  inv1  g1147(.a(n1027), .O(n1211));
  nand2 g1148(.a(n1062), .b(n1211), .O(n1212));
  nand2 g1149(.a(n1209), .b(n1211), .O(n1213));
  and2  g1150(.a(n1213), .b(n1212), .O(n1214));
  nand2 g1151(.a(n1214), .b(n1210), .O(n1215));
  xor2  g1152(.a(n1215), .b(n1208), .O(n1216));
  xor2  g1153(.a(n1216), .b(n1173), .O(n1217));
  nand2 g1154(.a(n1070), .b(n1063), .O(n1218));
  inv1  g1155(.a(n1026), .O(n1219));
  nand2 g1156(.a(n1070), .b(n1219), .O(n1220));
  nand2 g1157(.a(n1063), .b(n1219), .O(n1221));
  and2  g1158(.a(n1221), .b(n1220), .O(n1222));
  nand2 g1159(.a(n1222), .b(n1218), .O(n1223));
  xor2  g1160(.a(n1223), .b(n1217), .O(n1224));
  xor2  g1161(.a(n1224), .b(n1171), .O(n1225));
  inv1  g1162(.a(n1071), .O(n1226));
  nand2 g1163(.a(n1079), .b(n1226), .O(n1227));
  inv1  g1164(.a(n1025), .O(n1228));
  nand2 g1165(.a(n1079), .b(n1228), .O(n1229));
  nand2 g1166(.a(n1226), .b(n1228), .O(n1230));
  and2  g1167(.a(n1230), .b(n1229), .O(n1231));
  nand2 g1168(.a(n1231), .b(n1227), .O(n1232));
  xor2  g1169(.a(n1232), .b(n1225), .O(n1233));
  xor2  g1170(.a(n1233), .b(n1169), .O(n1234));
  nand2 g1171(.a(n1087), .b(n1080), .O(n1235));
  inv1  g1172(.a(n1024), .O(n1236));
  nand2 g1173(.a(n1087), .b(n1236), .O(n1237));
  nand2 g1174(.a(n1080), .b(n1236), .O(n1238));
  and2  g1175(.a(n1238), .b(n1237), .O(n1239));
  nand2 g1176(.a(n1239), .b(n1235), .O(n1240));
  xor2  g1177(.a(n1240), .b(n1234), .O(n1241));
  xor2  g1178(.a(n1241), .b(n1167), .O(n1242));
  inv1  g1179(.a(n1088), .O(n1243));
  nand2 g1180(.a(n1096), .b(n1243), .O(n1244));
  inv1  g1181(.a(n1023), .O(n1245));
  nand2 g1182(.a(n1096), .b(n1245), .O(n1246));
  nand2 g1183(.a(n1243), .b(n1245), .O(n1247));
  and2  g1184(.a(n1247), .b(n1246), .O(n1248));
  nand2 g1185(.a(n1248), .b(n1244), .O(n1249));
  xor2  g1186(.a(n1249), .b(n1242), .O(n1250));
  xor2  g1187(.a(n1250), .b(n1165), .O(n1251));
  nand2 g1188(.a(n1104), .b(n1097), .O(n1252));
  inv1  g1189(.a(n1022), .O(n1253));
  nand2 g1190(.a(n1104), .b(n1253), .O(n1254));
  nand2 g1191(.a(n1097), .b(n1253), .O(n1255));
  and2  g1192(.a(n1255), .b(n1254), .O(n1256));
  nand2 g1193(.a(n1256), .b(n1252), .O(n1257));
  xor2  g1194(.a(n1257), .b(n1251), .O(n1258));
  xor2  g1195(.a(n1258), .b(n1163), .O(n1259));
  inv1  g1196(.a(n1105), .O(n1260));
  nand2 g1197(.a(n1113), .b(n1260), .O(n1261));
  inv1  g1198(.a(n1021), .O(n1262));
  nand2 g1199(.a(n1113), .b(n1262), .O(n1263));
  nand2 g1200(.a(n1260), .b(n1262), .O(n1264));
  and2  g1201(.a(n1264), .b(n1263), .O(n1265));
  nand2 g1202(.a(n1265), .b(n1261), .O(n1266));
  xor2  g1203(.a(n1266), .b(n1259), .O(n1267));
  xor2  g1204(.a(n1267), .b(n1161), .O(n1268));
  nand2 g1205(.a(n1121), .b(n1114), .O(n1269));
  inv1  g1206(.a(n1020), .O(n1270));
  nand2 g1207(.a(n1121), .b(n1270), .O(n1271));
  nand2 g1208(.a(n1114), .b(n1270), .O(n1272));
  and2  g1209(.a(n1272), .b(n1271), .O(n1273));
  nand2 g1210(.a(n1273), .b(n1269), .O(n1274));
  xor2  g1211(.a(n1274), .b(n1268), .O(n1275));
  xor2  g1212(.a(n1275), .b(n1159), .O(n1276));
  inv1  g1213(.a(n1122), .O(n1277));
  nand2 g1214(.a(n1130), .b(n1277), .O(n1278));
  inv1  g1215(.a(n1019), .O(n1279));
  nand2 g1216(.a(n1130), .b(n1279), .O(n1280));
  nand2 g1217(.a(n1277), .b(n1279), .O(n1281));
  and2  g1218(.a(n1281), .b(n1280), .O(n1282));
  nand2 g1219(.a(n1282), .b(n1278), .O(n1283));
  xor2  g1220(.a(n1283), .b(n1276), .O(n1284));
  xor2  g1221(.a(n1284), .b(n1157), .O(n1285));
  nand2 g1222(.a(n1138), .b(n1131), .O(n1286));
  inv1  g1223(.a(n1018), .O(n1287));
  nand2 g1224(.a(n1138), .b(n1287), .O(n1288));
  nand2 g1225(.a(n1131), .b(n1287), .O(n1289));
  and2  g1226(.a(n1289), .b(n1288), .O(n1290));
  nand2 g1227(.a(n1290), .b(n1286), .O(n1291));
  xor2  g1228(.a(n1291), .b(n1285), .O(n1292));
  inv1  g1229(.a(n1292), .O(n1293));
  xor2  g1230(.a(n1293), .b(n1155), .O(n1294));
  inv1  g1231(.a(n1139), .O(n1295));
  nand2 g1232(.a(n1147), .b(n1295), .O(n1296));
  inv1  g1233(.a(n1017), .O(n1297));
  nand2 g1234(.a(n1147), .b(n1297), .O(n1298));
  nand2 g1235(.a(n1295), .b(n1297), .O(n1299));
  and2  g1236(.a(n1299), .b(n1298), .O(n1300));
  nand2 g1237(.a(n1300), .b(n1296), .O(n1301));
  xor2  g1238(.a(n1301), .b(n1294), .O(z17 ));
  nand2 g1239(.a(n1301), .b(n1155), .O(n1303));
  nand2 g1240(.a(n1301), .b(n1293), .O(n1304));
  nand2 g1241(.a(n1293), .b(n1155), .O(n1305));
  and2  g1242(.a(n1305), .b(n1304), .O(n1306));
  nand2 g1243(.a(n1306), .b(n1303), .O(n1307));
  nand2 g1244(.a(b15 ), .b(a3 ), .O(n1308));
  nand2 g1245(.a(b14 ), .b(a4 ), .O(n1309));
  inv1  g1246(.a(n1309), .O(n1310));
  nand2 g1247(.a(b13 ), .b(a5 ), .O(n1311));
  inv1  g1248(.a(n1311), .O(n1312));
  nand2 g1249(.a(b12 ), .b(a6 ), .O(n1313));
  inv1  g1250(.a(n1313), .O(n1314));
  nand2 g1251(.a(b11 ), .b(a7 ), .O(n1315));
  inv1  g1252(.a(n1315), .O(n1316));
  nand2 g1253(.a(b10 ), .b(a8 ), .O(n1317));
  inv1  g1254(.a(n1317), .O(n1318));
  nand2 g1255(.a(b9 ), .b(a9 ), .O(n1319));
  inv1  g1256(.a(n1319), .O(n1320));
  nand2 g1257(.a(b8 ), .b(a10 ), .O(n1321));
  inv1  g1258(.a(n1321), .O(n1322));
  nand2 g1259(.a(b7 ), .b(a11 ), .O(n1323));
  inv1  g1260(.a(n1323), .O(n1324));
  nand2 g1261(.a(b6 ), .b(a12 ), .O(n1325));
  inv1  g1262(.a(n1325), .O(n1326));
  nand2 g1263(.a(b5 ), .b(a13 ), .O(n1327));
  inv1  g1264(.a(n1327), .O(n1328));
  nand2 g1265(.a(b4 ), .b(a14 ), .O(n1329));
  nand2 g1266(.a(b3 ), .b(a15 ), .O(n1330));
  xnor2 g1267(.a(n1330), .b(n1329), .O(n1331));
  inv1  g1268(.a(n1181), .O(n1332));
  nand2 g1269(.a(n1190), .b(n1332), .O(n1333));
  inv1  g1270(.a(n1180), .O(n1334));
  nand2 g1271(.a(n1190), .b(n1334), .O(n1335));
  nand2 g1272(.a(n1332), .b(n1334), .O(n1336));
  and2  g1273(.a(n1336), .b(n1335), .O(n1337));
  nand2 g1274(.a(n1337), .b(n1333), .O(n1338));
  xor2  g1275(.a(n1338), .b(n1331), .O(n1339));
  xor2  g1276(.a(n1339), .b(n1328), .O(n1340));
  inv1  g1277(.a(n1191), .O(n1341));
  nand2 g1278(.a(n1198), .b(n1341), .O(n1342));
  nand2 g1279(.a(n1198), .b(n1179), .O(n1343));
  nand2 g1280(.a(n1341), .b(n1179), .O(n1344));
  and2  g1281(.a(n1344), .b(n1343), .O(n1345));
  nand2 g1282(.a(n1345), .b(n1342), .O(n1346));
  xor2  g1283(.a(n1346), .b(n1340), .O(n1347));
  xor2  g1284(.a(n1347), .b(n1326), .O(n1348));
  inv1  g1285(.a(n1199), .O(n1349));
  nand2 g1286(.a(n1206), .b(n1349), .O(n1350));
  nand2 g1287(.a(n1206), .b(n1177), .O(n1351));
  nand2 g1288(.a(n1349), .b(n1177), .O(n1352));
  and2  g1289(.a(n1352), .b(n1351), .O(n1353));
  nand2 g1290(.a(n1353), .b(n1350), .O(n1354));
  xor2  g1291(.a(n1354), .b(n1348), .O(n1355));
  xor2  g1292(.a(n1355), .b(n1324), .O(n1356));
  inv1  g1293(.a(n1207), .O(n1357));
  nand2 g1294(.a(n1215), .b(n1357), .O(n1358));
  nand2 g1295(.a(n1215), .b(n1175), .O(n1359));
  nand2 g1296(.a(n1357), .b(n1175), .O(n1360));
  and2  g1297(.a(n1360), .b(n1359), .O(n1361));
  nand2 g1298(.a(n1361), .b(n1358), .O(n1362));
  xor2  g1299(.a(n1362), .b(n1356), .O(n1363));
  xor2  g1300(.a(n1363), .b(n1322), .O(n1364));
  inv1  g1301(.a(n1216), .O(n1365));
  nand2 g1302(.a(n1223), .b(n1365), .O(n1366));
  nand2 g1303(.a(n1223), .b(n1173), .O(n1367));
  nand2 g1304(.a(n1365), .b(n1173), .O(n1368));
  and2  g1305(.a(n1368), .b(n1367), .O(n1369));
  nand2 g1306(.a(n1369), .b(n1366), .O(n1370));
  xor2  g1307(.a(n1370), .b(n1364), .O(n1371));
  xor2  g1308(.a(n1371), .b(n1320), .O(n1372));
  inv1  g1309(.a(n1224), .O(n1373));
  nand2 g1310(.a(n1232), .b(n1373), .O(n1374));
  nand2 g1311(.a(n1232), .b(n1171), .O(n1375));
  nand2 g1312(.a(n1373), .b(n1171), .O(n1376));
  and2  g1313(.a(n1376), .b(n1375), .O(n1377));
  nand2 g1314(.a(n1377), .b(n1374), .O(n1378));
  xor2  g1315(.a(n1378), .b(n1372), .O(n1379));
  xor2  g1316(.a(n1379), .b(n1318), .O(n1380));
  inv1  g1317(.a(n1233), .O(n1381));
  nand2 g1318(.a(n1240), .b(n1381), .O(n1382));
  nand2 g1319(.a(n1240), .b(n1169), .O(n1383));
  nand2 g1320(.a(n1381), .b(n1169), .O(n1384));
  and2  g1321(.a(n1384), .b(n1383), .O(n1385));
  nand2 g1322(.a(n1385), .b(n1382), .O(n1386));
  xor2  g1323(.a(n1386), .b(n1380), .O(n1387));
  xor2  g1324(.a(n1387), .b(n1316), .O(n1388));
  inv1  g1325(.a(n1241), .O(n1389));
  nand2 g1326(.a(n1249), .b(n1389), .O(n1390));
  nand2 g1327(.a(n1249), .b(n1167), .O(n1391));
  nand2 g1328(.a(n1389), .b(n1167), .O(n1392));
  and2  g1329(.a(n1392), .b(n1391), .O(n1393));
  nand2 g1330(.a(n1393), .b(n1390), .O(n1394));
  xor2  g1331(.a(n1394), .b(n1388), .O(n1395));
  xor2  g1332(.a(n1395), .b(n1314), .O(n1396));
  inv1  g1333(.a(n1250), .O(n1397));
  nand2 g1334(.a(n1257), .b(n1397), .O(n1398));
  nand2 g1335(.a(n1257), .b(n1165), .O(n1399));
  nand2 g1336(.a(n1397), .b(n1165), .O(n1400));
  and2  g1337(.a(n1400), .b(n1399), .O(n1401));
  nand2 g1338(.a(n1401), .b(n1398), .O(n1402));
  xor2  g1339(.a(n1402), .b(n1396), .O(n1403));
  xor2  g1340(.a(n1403), .b(n1312), .O(n1404));
  inv1  g1341(.a(n1258), .O(n1405));
  nand2 g1342(.a(n1266), .b(n1405), .O(n1406));
  nand2 g1343(.a(n1266), .b(n1163), .O(n1407));
  nand2 g1344(.a(n1405), .b(n1163), .O(n1408));
  and2  g1345(.a(n1408), .b(n1407), .O(n1409));
  nand2 g1346(.a(n1409), .b(n1406), .O(n1410));
  xor2  g1347(.a(n1410), .b(n1404), .O(n1411));
  xor2  g1348(.a(n1411), .b(n1310), .O(n1412));
  inv1  g1349(.a(n1267), .O(n1413));
  nand2 g1350(.a(n1274), .b(n1413), .O(n1414));
  nand2 g1351(.a(n1274), .b(n1161), .O(n1415));
  nand2 g1352(.a(n1413), .b(n1161), .O(n1416));
  and2  g1353(.a(n1416), .b(n1415), .O(n1417));
  nand2 g1354(.a(n1417), .b(n1414), .O(n1418));
  xor2  g1355(.a(n1418), .b(n1412), .O(n1419));
  xor2  g1356(.a(n1419), .b(n1308), .O(n1420));
  inv1  g1357(.a(n1275), .O(n1421));
  nand2 g1358(.a(n1283), .b(n1421), .O(n1422));
  nand2 g1359(.a(n1283), .b(n1159), .O(n1423));
  nand2 g1360(.a(n1421), .b(n1159), .O(n1424));
  and2  g1361(.a(n1424), .b(n1423), .O(n1425));
  nand2 g1362(.a(n1425), .b(n1422), .O(n1426));
  xor2  g1363(.a(n1426), .b(n1420), .O(n1427));
  xor2  g1364(.a(n1427), .b(n1307), .O(n1428));
  inv1  g1365(.a(n1284), .O(n1429));
  nand2 g1366(.a(n1291), .b(n1429), .O(n1430));
  nand2 g1367(.a(n1291), .b(n1157), .O(n1431));
  nand2 g1368(.a(n1429), .b(n1157), .O(n1432));
  and2  g1369(.a(n1432), .b(n1431), .O(n1433));
  nand2 g1370(.a(n1433), .b(n1430), .O(n1434));
  xor2  g1371(.a(n1434), .b(n1428), .O(z18 ));
  nand2 g1372(.a(n1434), .b(n1307), .O(n1436));
  nand2 g1373(.a(n1434), .b(n1427), .O(n1437));
  nand2 g1374(.a(n1427), .b(n1307), .O(n1438));
  and2  g1375(.a(n1438), .b(n1437), .O(n1439));
  nand2 g1376(.a(n1439), .b(n1436), .O(n1440));
  nand2 g1377(.a(b15 ), .b(a4 ), .O(n1441));
  nand2 g1378(.a(b14 ), .b(a5 ), .O(n1442));
  inv1  g1379(.a(n1442), .O(n1443));
  nand2 g1380(.a(b13 ), .b(a6 ), .O(n1444));
  inv1  g1381(.a(n1444), .O(n1445));
  nand2 g1382(.a(b12 ), .b(a7 ), .O(n1446));
  inv1  g1383(.a(n1446), .O(n1447));
  nand2 g1384(.a(b11 ), .b(a8 ), .O(n1448));
  inv1  g1385(.a(n1448), .O(n1449));
  nand2 g1386(.a(b10 ), .b(a9 ), .O(n1450));
  inv1  g1387(.a(n1450), .O(n1451));
  nand2 g1388(.a(b9 ), .b(a10 ), .O(n1452));
  inv1  g1389(.a(n1452), .O(n1453));
  nand2 g1390(.a(b8 ), .b(a11 ), .O(n1454));
  inv1  g1391(.a(n1454), .O(n1455));
  nand2 g1392(.a(b7 ), .b(a12 ), .O(n1456));
  inv1  g1393(.a(n1456), .O(n1457));
  nand2 g1394(.a(b6 ), .b(a13 ), .O(n1458));
  inv1  g1395(.a(n1458), .O(n1459));
  nand2 g1396(.a(b5 ), .b(a14 ), .O(n1460));
  nand2 g1397(.a(b4 ), .b(a15 ), .O(n1461));
  xnor2 g1398(.a(n1461), .b(n1460), .O(n1462));
  inv1  g1399(.a(n1330), .O(n1463));
  nand2 g1400(.a(n1338), .b(n1463), .O(n1464));
  inv1  g1401(.a(n1329), .O(n1465));
  nand2 g1402(.a(n1338), .b(n1465), .O(n1466));
  nand2 g1403(.a(n1463), .b(n1465), .O(n1467));
  and2  g1404(.a(n1467), .b(n1466), .O(n1468));
  nand2 g1405(.a(n1468), .b(n1464), .O(n1469));
  xor2  g1406(.a(n1469), .b(n1462), .O(n1470));
  xor2  g1407(.a(n1470), .b(n1459), .O(n1471));
  inv1  g1408(.a(n1339), .O(n1472));
  nand2 g1409(.a(n1346), .b(n1472), .O(n1473));
  nand2 g1410(.a(n1346), .b(n1328), .O(n1474));
  nand2 g1411(.a(n1472), .b(n1328), .O(n1475));
  and2  g1412(.a(n1475), .b(n1474), .O(n1476));
  nand2 g1413(.a(n1476), .b(n1473), .O(n1477));
  xor2  g1414(.a(n1477), .b(n1471), .O(n1478));
  xor2  g1415(.a(n1478), .b(n1457), .O(n1479));
  inv1  g1416(.a(n1347), .O(n1480));
  nand2 g1417(.a(n1354), .b(n1480), .O(n1481));
  nand2 g1418(.a(n1354), .b(n1326), .O(n1482));
  nand2 g1419(.a(n1480), .b(n1326), .O(n1483));
  and2  g1420(.a(n1483), .b(n1482), .O(n1484));
  nand2 g1421(.a(n1484), .b(n1481), .O(n1485));
  xor2  g1422(.a(n1485), .b(n1479), .O(n1486));
  xor2  g1423(.a(n1486), .b(n1455), .O(n1487));
  inv1  g1424(.a(n1355), .O(n1488));
  nand2 g1425(.a(n1362), .b(n1488), .O(n1489));
  nand2 g1426(.a(n1362), .b(n1324), .O(n1490));
  nand2 g1427(.a(n1488), .b(n1324), .O(n1491));
  and2  g1428(.a(n1491), .b(n1490), .O(n1492));
  nand2 g1429(.a(n1492), .b(n1489), .O(n1493));
  xor2  g1430(.a(n1493), .b(n1487), .O(n1494));
  xor2  g1431(.a(n1494), .b(n1453), .O(n1495));
  inv1  g1432(.a(n1363), .O(n1496));
  nand2 g1433(.a(n1370), .b(n1496), .O(n1497));
  nand2 g1434(.a(n1370), .b(n1322), .O(n1498));
  nand2 g1435(.a(n1496), .b(n1322), .O(n1499));
  and2  g1436(.a(n1499), .b(n1498), .O(n1500));
  nand2 g1437(.a(n1500), .b(n1497), .O(n1501));
  xor2  g1438(.a(n1501), .b(n1495), .O(n1502));
  xor2  g1439(.a(n1502), .b(n1451), .O(n1503));
  inv1  g1440(.a(n1371), .O(n1504));
  nand2 g1441(.a(n1378), .b(n1504), .O(n1505));
  nand2 g1442(.a(n1378), .b(n1320), .O(n1506));
  nand2 g1443(.a(n1504), .b(n1320), .O(n1507));
  and2  g1444(.a(n1507), .b(n1506), .O(n1508));
  nand2 g1445(.a(n1508), .b(n1505), .O(n1509));
  xor2  g1446(.a(n1509), .b(n1503), .O(n1510));
  xor2  g1447(.a(n1510), .b(n1449), .O(n1511));
  inv1  g1448(.a(n1379), .O(n1512));
  nand2 g1449(.a(n1386), .b(n1512), .O(n1513));
  nand2 g1450(.a(n1386), .b(n1318), .O(n1514));
  nand2 g1451(.a(n1512), .b(n1318), .O(n1515));
  and2  g1452(.a(n1515), .b(n1514), .O(n1516));
  nand2 g1453(.a(n1516), .b(n1513), .O(n1517));
  xor2  g1454(.a(n1517), .b(n1511), .O(n1518));
  xor2  g1455(.a(n1518), .b(n1447), .O(n1519));
  inv1  g1456(.a(n1387), .O(n1520));
  nand2 g1457(.a(n1394), .b(n1520), .O(n1521));
  nand2 g1458(.a(n1394), .b(n1316), .O(n1522));
  nand2 g1459(.a(n1520), .b(n1316), .O(n1523));
  and2  g1460(.a(n1523), .b(n1522), .O(n1524));
  nand2 g1461(.a(n1524), .b(n1521), .O(n1525));
  xor2  g1462(.a(n1525), .b(n1519), .O(n1526));
  xor2  g1463(.a(n1526), .b(n1445), .O(n1527));
  inv1  g1464(.a(n1395), .O(n1528));
  nand2 g1465(.a(n1402), .b(n1528), .O(n1529));
  nand2 g1466(.a(n1402), .b(n1314), .O(n1530));
  nand2 g1467(.a(n1528), .b(n1314), .O(n1531));
  and2  g1468(.a(n1531), .b(n1530), .O(n1532));
  nand2 g1469(.a(n1532), .b(n1529), .O(n1533));
  xor2  g1470(.a(n1533), .b(n1527), .O(n1534));
  xor2  g1471(.a(n1534), .b(n1443), .O(n1535));
  inv1  g1472(.a(n1403), .O(n1536));
  nand2 g1473(.a(n1410), .b(n1536), .O(n1537));
  nand2 g1474(.a(n1410), .b(n1312), .O(n1538));
  nand2 g1475(.a(n1536), .b(n1312), .O(n1539));
  and2  g1476(.a(n1539), .b(n1538), .O(n1540));
  nand2 g1477(.a(n1540), .b(n1537), .O(n1541));
  xor2  g1478(.a(n1541), .b(n1535), .O(n1542));
  xor2  g1479(.a(n1542), .b(n1441), .O(n1543));
  inv1  g1480(.a(n1411), .O(n1544));
  nand2 g1481(.a(n1418), .b(n1544), .O(n1545));
  nand2 g1482(.a(n1418), .b(n1310), .O(n1546));
  nand2 g1483(.a(n1544), .b(n1310), .O(n1547));
  and2  g1484(.a(n1547), .b(n1546), .O(n1548));
  nand2 g1485(.a(n1548), .b(n1545), .O(n1549));
  xor2  g1486(.a(n1549), .b(n1543), .O(n1550));
  xor2  g1487(.a(n1550), .b(n1440), .O(n1551));
  inv1  g1488(.a(n1419), .O(n1552));
  nand2 g1489(.a(n1426), .b(n1552), .O(n1553));
  inv1  g1490(.a(n1308), .O(n1554));
  nand2 g1491(.a(n1426), .b(n1554), .O(n1555));
  nand2 g1492(.a(n1552), .b(n1554), .O(n1556));
  and2  g1493(.a(n1556), .b(n1555), .O(n1557));
  nand2 g1494(.a(n1557), .b(n1553), .O(n1558));
  xor2  g1495(.a(n1558), .b(n1551), .O(z19 ));
  nand2 g1496(.a(n1558), .b(n1440), .O(n1560));
  nand2 g1497(.a(n1558), .b(n1550), .O(n1561));
  nand2 g1498(.a(n1550), .b(n1440), .O(n1562));
  and2  g1499(.a(n1562), .b(n1561), .O(n1563));
  nand2 g1500(.a(n1563), .b(n1560), .O(n1564));
  nand2 g1501(.a(b15 ), .b(a5 ), .O(n1565));
  nand2 g1502(.a(b14 ), .b(a6 ), .O(n1566));
  inv1  g1503(.a(n1566), .O(n1567));
  nand2 g1504(.a(b13 ), .b(a7 ), .O(n1568));
  inv1  g1505(.a(n1568), .O(n1569));
  nand2 g1506(.a(b12 ), .b(a8 ), .O(n1570));
  inv1  g1507(.a(n1570), .O(n1571));
  nand2 g1508(.a(b11 ), .b(a9 ), .O(n1572));
  inv1  g1509(.a(n1572), .O(n1573));
  nand2 g1510(.a(b10 ), .b(a10 ), .O(n1574));
  inv1  g1511(.a(n1574), .O(n1575));
  nand2 g1512(.a(b9 ), .b(a11 ), .O(n1576));
  inv1  g1513(.a(n1576), .O(n1577));
  nand2 g1514(.a(b8 ), .b(a12 ), .O(n1578));
  inv1  g1515(.a(n1578), .O(n1579));
  nand2 g1516(.a(b7 ), .b(a13 ), .O(n1580));
  inv1  g1517(.a(n1580), .O(n1581));
  nand2 g1518(.a(b6 ), .b(a14 ), .O(n1582));
  nand2 g1519(.a(b5 ), .b(a15 ), .O(n1583));
  xnor2 g1520(.a(n1583), .b(n1582), .O(n1584));
  inv1  g1521(.a(n1461), .O(n1585));
  nand2 g1522(.a(n1469), .b(n1585), .O(n1586));
  inv1  g1523(.a(n1460), .O(n1587));
  nand2 g1524(.a(n1469), .b(n1587), .O(n1588));
  nand2 g1525(.a(n1585), .b(n1587), .O(n1589));
  and2  g1526(.a(n1589), .b(n1588), .O(n1590));
  nand2 g1527(.a(n1590), .b(n1586), .O(n1591));
  xor2  g1528(.a(n1591), .b(n1584), .O(n1592));
  xor2  g1529(.a(n1592), .b(n1581), .O(n1593));
  inv1  g1530(.a(n1470), .O(n1594));
  nand2 g1531(.a(n1477), .b(n1594), .O(n1595));
  nand2 g1532(.a(n1477), .b(n1459), .O(n1596));
  nand2 g1533(.a(n1594), .b(n1459), .O(n1597));
  and2  g1534(.a(n1597), .b(n1596), .O(n1598));
  nand2 g1535(.a(n1598), .b(n1595), .O(n1599));
  xor2  g1536(.a(n1599), .b(n1593), .O(n1600));
  xor2  g1537(.a(n1600), .b(n1579), .O(n1601));
  inv1  g1538(.a(n1478), .O(n1602));
  nand2 g1539(.a(n1485), .b(n1602), .O(n1603));
  nand2 g1540(.a(n1485), .b(n1457), .O(n1604));
  nand2 g1541(.a(n1602), .b(n1457), .O(n1605));
  and2  g1542(.a(n1605), .b(n1604), .O(n1606));
  nand2 g1543(.a(n1606), .b(n1603), .O(n1607));
  xor2  g1544(.a(n1607), .b(n1601), .O(n1608));
  xor2  g1545(.a(n1608), .b(n1577), .O(n1609));
  inv1  g1546(.a(n1486), .O(n1610));
  nand2 g1547(.a(n1493), .b(n1610), .O(n1611));
  nand2 g1548(.a(n1493), .b(n1455), .O(n1612));
  nand2 g1549(.a(n1610), .b(n1455), .O(n1613));
  and2  g1550(.a(n1613), .b(n1612), .O(n1614));
  nand2 g1551(.a(n1614), .b(n1611), .O(n1615));
  xor2  g1552(.a(n1615), .b(n1609), .O(n1616));
  xor2  g1553(.a(n1616), .b(n1575), .O(n1617));
  inv1  g1554(.a(n1494), .O(n1618));
  nand2 g1555(.a(n1501), .b(n1618), .O(n1619));
  nand2 g1556(.a(n1501), .b(n1453), .O(n1620));
  nand2 g1557(.a(n1618), .b(n1453), .O(n1621));
  and2  g1558(.a(n1621), .b(n1620), .O(n1622));
  nand2 g1559(.a(n1622), .b(n1619), .O(n1623));
  xor2  g1560(.a(n1623), .b(n1617), .O(n1624));
  xor2  g1561(.a(n1624), .b(n1573), .O(n1625));
  inv1  g1562(.a(n1502), .O(n1626));
  nand2 g1563(.a(n1509), .b(n1626), .O(n1627));
  nand2 g1564(.a(n1509), .b(n1451), .O(n1628));
  nand2 g1565(.a(n1626), .b(n1451), .O(n1629));
  and2  g1566(.a(n1629), .b(n1628), .O(n1630));
  nand2 g1567(.a(n1630), .b(n1627), .O(n1631));
  xor2  g1568(.a(n1631), .b(n1625), .O(n1632));
  xor2  g1569(.a(n1632), .b(n1571), .O(n1633));
  inv1  g1570(.a(n1510), .O(n1634));
  nand2 g1571(.a(n1517), .b(n1634), .O(n1635));
  nand2 g1572(.a(n1517), .b(n1449), .O(n1636));
  nand2 g1573(.a(n1634), .b(n1449), .O(n1637));
  and2  g1574(.a(n1637), .b(n1636), .O(n1638));
  nand2 g1575(.a(n1638), .b(n1635), .O(n1639));
  xor2  g1576(.a(n1639), .b(n1633), .O(n1640));
  xor2  g1577(.a(n1640), .b(n1569), .O(n1641));
  inv1  g1578(.a(n1518), .O(n1642));
  nand2 g1579(.a(n1525), .b(n1642), .O(n1643));
  nand2 g1580(.a(n1525), .b(n1447), .O(n1644));
  nand2 g1581(.a(n1642), .b(n1447), .O(n1645));
  and2  g1582(.a(n1645), .b(n1644), .O(n1646));
  nand2 g1583(.a(n1646), .b(n1643), .O(n1647));
  xor2  g1584(.a(n1647), .b(n1641), .O(n1648));
  xor2  g1585(.a(n1648), .b(n1567), .O(n1649));
  inv1  g1586(.a(n1526), .O(n1650));
  nand2 g1587(.a(n1533), .b(n1650), .O(n1651));
  nand2 g1588(.a(n1533), .b(n1445), .O(n1652));
  nand2 g1589(.a(n1650), .b(n1445), .O(n1653));
  and2  g1590(.a(n1653), .b(n1652), .O(n1654));
  nand2 g1591(.a(n1654), .b(n1651), .O(n1655));
  xor2  g1592(.a(n1655), .b(n1649), .O(n1656));
  xor2  g1593(.a(n1656), .b(n1565), .O(n1657));
  inv1  g1594(.a(n1534), .O(n1658));
  nand2 g1595(.a(n1541), .b(n1658), .O(n1659));
  nand2 g1596(.a(n1541), .b(n1443), .O(n1660));
  nand2 g1597(.a(n1658), .b(n1443), .O(n1661));
  and2  g1598(.a(n1661), .b(n1660), .O(n1662));
  nand2 g1599(.a(n1662), .b(n1659), .O(n1663));
  xor2  g1600(.a(n1663), .b(n1657), .O(n1664));
  xor2  g1601(.a(n1664), .b(n1564), .O(n1665));
  inv1  g1602(.a(n1542), .O(n1666));
  nand2 g1603(.a(n1549), .b(n1666), .O(n1667));
  inv1  g1604(.a(n1441), .O(n1668));
  nand2 g1605(.a(n1549), .b(n1668), .O(n1669));
  nand2 g1606(.a(n1666), .b(n1668), .O(n1670));
  and2  g1607(.a(n1670), .b(n1669), .O(n1671));
  nand2 g1608(.a(n1671), .b(n1667), .O(n1672));
  xor2  g1609(.a(n1672), .b(n1665), .O(z20 ));
  nand2 g1610(.a(n1672), .b(n1564), .O(n1674));
  nand2 g1611(.a(n1672), .b(n1664), .O(n1675));
  nand2 g1612(.a(n1664), .b(n1564), .O(n1676));
  and2  g1613(.a(n1676), .b(n1675), .O(n1677));
  nand2 g1614(.a(n1677), .b(n1674), .O(n1678));
  nand2 g1615(.a(b15 ), .b(a6 ), .O(n1679));
  nand2 g1616(.a(b14 ), .b(a7 ), .O(n1680));
  inv1  g1617(.a(n1680), .O(n1681));
  nand2 g1618(.a(b13 ), .b(a8 ), .O(n1682));
  inv1  g1619(.a(n1682), .O(n1683));
  nand2 g1620(.a(b12 ), .b(a9 ), .O(n1684));
  inv1  g1621(.a(n1684), .O(n1685));
  nand2 g1622(.a(b11 ), .b(a10 ), .O(n1686));
  inv1  g1623(.a(n1686), .O(n1687));
  nand2 g1624(.a(b10 ), .b(a11 ), .O(n1688));
  inv1  g1625(.a(n1688), .O(n1689));
  nand2 g1626(.a(b9 ), .b(a12 ), .O(n1690));
  inv1  g1627(.a(n1690), .O(n1691));
  nand2 g1628(.a(b8 ), .b(a13 ), .O(n1692));
  inv1  g1629(.a(n1692), .O(n1693));
  nand2 g1630(.a(b7 ), .b(a14 ), .O(n1694));
  nand2 g1631(.a(b6 ), .b(a15 ), .O(n1695));
  xnor2 g1632(.a(n1695), .b(n1694), .O(n1696));
  inv1  g1633(.a(n1583), .O(n1697));
  nand2 g1634(.a(n1591), .b(n1697), .O(n1698));
  inv1  g1635(.a(n1582), .O(n1699));
  nand2 g1636(.a(n1591), .b(n1699), .O(n1700));
  nand2 g1637(.a(n1697), .b(n1699), .O(n1701));
  and2  g1638(.a(n1701), .b(n1700), .O(n1702));
  nand2 g1639(.a(n1702), .b(n1698), .O(n1703));
  xor2  g1640(.a(n1703), .b(n1696), .O(n1704));
  xor2  g1641(.a(n1704), .b(n1693), .O(n1705));
  inv1  g1642(.a(n1592), .O(n1706));
  nand2 g1643(.a(n1599), .b(n1706), .O(n1707));
  nand2 g1644(.a(n1599), .b(n1581), .O(n1708));
  nand2 g1645(.a(n1706), .b(n1581), .O(n1709));
  and2  g1646(.a(n1709), .b(n1708), .O(n1710));
  nand2 g1647(.a(n1710), .b(n1707), .O(n1711));
  xor2  g1648(.a(n1711), .b(n1705), .O(n1712));
  xor2  g1649(.a(n1712), .b(n1691), .O(n1713));
  inv1  g1650(.a(n1600), .O(n1714));
  nand2 g1651(.a(n1607), .b(n1714), .O(n1715));
  nand2 g1652(.a(n1607), .b(n1579), .O(n1716));
  nand2 g1653(.a(n1714), .b(n1579), .O(n1717));
  and2  g1654(.a(n1717), .b(n1716), .O(n1718));
  nand2 g1655(.a(n1718), .b(n1715), .O(n1719));
  xor2  g1656(.a(n1719), .b(n1713), .O(n1720));
  xor2  g1657(.a(n1720), .b(n1689), .O(n1721));
  inv1  g1658(.a(n1608), .O(n1722));
  nand2 g1659(.a(n1615), .b(n1722), .O(n1723));
  nand2 g1660(.a(n1615), .b(n1577), .O(n1724));
  nand2 g1661(.a(n1722), .b(n1577), .O(n1725));
  and2  g1662(.a(n1725), .b(n1724), .O(n1726));
  nand2 g1663(.a(n1726), .b(n1723), .O(n1727));
  xor2  g1664(.a(n1727), .b(n1721), .O(n1728));
  xor2  g1665(.a(n1728), .b(n1687), .O(n1729));
  inv1  g1666(.a(n1616), .O(n1730));
  nand2 g1667(.a(n1623), .b(n1730), .O(n1731));
  nand2 g1668(.a(n1623), .b(n1575), .O(n1732));
  nand2 g1669(.a(n1730), .b(n1575), .O(n1733));
  and2  g1670(.a(n1733), .b(n1732), .O(n1734));
  nand2 g1671(.a(n1734), .b(n1731), .O(n1735));
  xor2  g1672(.a(n1735), .b(n1729), .O(n1736));
  xor2  g1673(.a(n1736), .b(n1685), .O(n1737));
  inv1  g1674(.a(n1624), .O(n1738));
  nand2 g1675(.a(n1631), .b(n1738), .O(n1739));
  nand2 g1676(.a(n1631), .b(n1573), .O(n1740));
  nand2 g1677(.a(n1738), .b(n1573), .O(n1741));
  and2  g1678(.a(n1741), .b(n1740), .O(n1742));
  nand2 g1679(.a(n1742), .b(n1739), .O(n1743));
  xor2  g1680(.a(n1743), .b(n1737), .O(n1744));
  xor2  g1681(.a(n1744), .b(n1683), .O(n1745));
  inv1  g1682(.a(n1632), .O(n1746));
  nand2 g1683(.a(n1639), .b(n1746), .O(n1747));
  nand2 g1684(.a(n1639), .b(n1571), .O(n1748));
  nand2 g1685(.a(n1746), .b(n1571), .O(n1749));
  and2  g1686(.a(n1749), .b(n1748), .O(n1750));
  nand2 g1687(.a(n1750), .b(n1747), .O(n1751));
  xor2  g1688(.a(n1751), .b(n1745), .O(n1752));
  xor2  g1689(.a(n1752), .b(n1681), .O(n1753));
  inv1  g1690(.a(n1640), .O(n1754));
  nand2 g1691(.a(n1647), .b(n1754), .O(n1755));
  nand2 g1692(.a(n1647), .b(n1569), .O(n1756));
  nand2 g1693(.a(n1754), .b(n1569), .O(n1757));
  and2  g1694(.a(n1757), .b(n1756), .O(n1758));
  nand2 g1695(.a(n1758), .b(n1755), .O(n1759));
  xor2  g1696(.a(n1759), .b(n1753), .O(n1760));
  xor2  g1697(.a(n1760), .b(n1679), .O(n1761));
  inv1  g1698(.a(n1648), .O(n1762));
  nand2 g1699(.a(n1655), .b(n1762), .O(n1763));
  nand2 g1700(.a(n1655), .b(n1567), .O(n1764));
  nand2 g1701(.a(n1762), .b(n1567), .O(n1765));
  and2  g1702(.a(n1765), .b(n1764), .O(n1766));
  nand2 g1703(.a(n1766), .b(n1763), .O(n1767));
  xor2  g1704(.a(n1767), .b(n1761), .O(n1768));
  xor2  g1705(.a(n1768), .b(n1678), .O(n1769));
  inv1  g1706(.a(n1656), .O(n1770));
  nand2 g1707(.a(n1663), .b(n1770), .O(n1771));
  inv1  g1708(.a(n1565), .O(n1772));
  nand2 g1709(.a(n1663), .b(n1772), .O(n1773));
  nand2 g1710(.a(n1770), .b(n1772), .O(n1774));
  and2  g1711(.a(n1774), .b(n1773), .O(n1775));
  nand2 g1712(.a(n1775), .b(n1771), .O(n1776));
  xor2  g1713(.a(n1776), .b(n1769), .O(z21 ));
  nand2 g1714(.a(n1776), .b(n1678), .O(n1778));
  nand2 g1715(.a(n1776), .b(n1768), .O(n1779));
  nand2 g1716(.a(n1768), .b(n1678), .O(n1780));
  and2  g1717(.a(n1780), .b(n1779), .O(n1781));
  nand2 g1718(.a(n1781), .b(n1778), .O(n1782));
  nand2 g1719(.a(b15 ), .b(a7 ), .O(n1783));
  nand2 g1720(.a(b14 ), .b(a8 ), .O(n1784));
  inv1  g1721(.a(n1784), .O(n1785));
  nand2 g1722(.a(b13 ), .b(a9 ), .O(n1786));
  inv1  g1723(.a(n1786), .O(n1787));
  nand2 g1724(.a(b12 ), .b(a10 ), .O(n1788));
  inv1  g1725(.a(n1788), .O(n1789));
  nand2 g1726(.a(b11 ), .b(a11 ), .O(n1790));
  inv1  g1727(.a(n1790), .O(n1791));
  nand2 g1728(.a(b10 ), .b(a12 ), .O(n1792));
  inv1  g1729(.a(n1792), .O(n1793));
  nand2 g1730(.a(b9 ), .b(a13 ), .O(n1794));
  inv1  g1731(.a(n1794), .O(n1795));
  nand2 g1732(.a(b8 ), .b(a14 ), .O(n1796));
  nand2 g1733(.a(b7 ), .b(a15 ), .O(n1797));
  xnor2 g1734(.a(n1797), .b(n1796), .O(n1798));
  inv1  g1735(.a(n1695), .O(n1799));
  nand2 g1736(.a(n1703), .b(n1799), .O(n1800));
  inv1  g1737(.a(n1694), .O(n1801));
  nand2 g1738(.a(n1703), .b(n1801), .O(n1802));
  nand2 g1739(.a(n1799), .b(n1801), .O(n1803));
  and2  g1740(.a(n1803), .b(n1802), .O(n1804));
  nand2 g1741(.a(n1804), .b(n1800), .O(n1805));
  xor2  g1742(.a(n1805), .b(n1798), .O(n1806));
  xor2  g1743(.a(n1806), .b(n1795), .O(n1807));
  inv1  g1744(.a(n1704), .O(n1808));
  nand2 g1745(.a(n1711), .b(n1808), .O(n1809));
  nand2 g1746(.a(n1711), .b(n1693), .O(n1810));
  nand2 g1747(.a(n1808), .b(n1693), .O(n1811));
  and2  g1748(.a(n1811), .b(n1810), .O(n1812));
  nand2 g1749(.a(n1812), .b(n1809), .O(n1813));
  xor2  g1750(.a(n1813), .b(n1807), .O(n1814));
  xor2  g1751(.a(n1814), .b(n1793), .O(n1815));
  inv1  g1752(.a(n1712), .O(n1816));
  nand2 g1753(.a(n1719), .b(n1816), .O(n1817));
  nand2 g1754(.a(n1719), .b(n1691), .O(n1818));
  nand2 g1755(.a(n1816), .b(n1691), .O(n1819));
  and2  g1756(.a(n1819), .b(n1818), .O(n1820));
  nand2 g1757(.a(n1820), .b(n1817), .O(n1821));
  xor2  g1758(.a(n1821), .b(n1815), .O(n1822));
  xor2  g1759(.a(n1822), .b(n1791), .O(n1823));
  inv1  g1760(.a(n1720), .O(n1824));
  nand2 g1761(.a(n1727), .b(n1824), .O(n1825));
  nand2 g1762(.a(n1727), .b(n1689), .O(n1826));
  nand2 g1763(.a(n1824), .b(n1689), .O(n1827));
  and2  g1764(.a(n1827), .b(n1826), .O(n1828));
  nand2 g1765(.a(n1828), .b(n1825), .O(n1829));
  xor2  g1766(.a(n1829), .b(n1823), .O(n1830));
  xor2  g1767(.a(n1830), .b(n1789), .O(n1831));
  inv1  g1768(.a(n1728), .O(n1832));
  nand2 g1769(.a(n1735), .b(n1832), .O(n1833));
  nand2 g1770(.a(n1735), .b(n1687), .O(n1834));
  nand2 g1771(.a(n1832), .b(n1687), .O(n1835));
  and2  g1772(.a(n1835), .b(n1834), .O(n1836));
  nand2 g1773(.a(n1836), .b(n1833), .O(n1837));
  xor2  g1774(.a(n1837), .b(n1831), .O(n1838));
  xor2  g1775(.a(n1838), .b(n1787), .O(n1839));
  inv1  g1776(.a(n1736), .O(n1840));
  nand2 g1777(.a(n1743), .b(n1840), .O(n1841));
  nand2 g1778(.a(n1743), .b(n1685), .O(n1842));
  nand2 g1779(.a(n1840), .b(n1685), .O(n1843));
  and2  g1780(.a(n1843), .b(n1842), .O(n1844));
  nand2 g1781(.a(n1844), .b(n1841), .O(n1845));
  xor2  g1782(.a(n1845), .b(n1839), .O(n1846));
  xor2  g1783(.a(n1846), .b(n1785), .O(n1847));
  inv1  g1784(.a(n1744), .O(n1848));
  nand2 g1785(.a(n1751), .b(n1848), .O(n1849));
  nand2 g1786(.a(n1751), .b(n1683), .O(n1850));
  nand2 g1787(.a(n1848), .b(n1683), .O(n1851));
  and2  g1788(.a(n1851), .b(n1850), .O(n1852));
  nand2 g1789(.a(n1852), .b(n1849), .O(n1853));
  xor2  g1790(.a(n1853), .b(n1847), .O(n1854));
  xor2  g1791(.a(n1854), .b(n1783), .O(n1855));
  inv1  g1792(.a(n1752), .O(n1856));
  nand2 g1793(.a(n1759), .b(n1856), .O(n1857));
  nand2 g1794(.a(n1759), .b(n1681), .O(n1858));
  nand2 g1795(.a(n1856), .b(n1681), .O(n1859));
  and2  g1796(.a(n1859), .b(n1858), .O(n1860));
  nand2 g1797(.a(n1860), .b(n1857), .O(n1861));
  xor2  g1798(.a(n1861), .b(n1855), .O(n1862));
  xor2  g1799(.a(n1862), .b(n1782), .O(n1863));
  inv1  g1800(.a(n1760), .O(n1864));
  nand2 g1801(.a(n1767), .b(n1864), .O(n1865));
  inv1  g1802(.a(n1679), .O(n1866));
  nand2 g1803(.a(n1767), .b(n1866), .O(n1867));
  nand2 g1804(.a(n1864), .b(n1866), .O(n1868));
  and2  g1805(.a(n1868), .b(n1867), .O(n1869));
  nand2 g1806(.a(n1869), .b(n1865), .O(n1870));
  xor2  g1807(.a(n1870), .b(n1863), .O(z22 ));
  nand2 g1808(.a(n1870), .b(n1782), .O(n1872));
  nand2 g1809(.a(n1870), .b(n1862), .O(n1873));
  nand2 g1810(.a(n1862), .b(n1782), .O(n1874));
  and2  g1811(.a(n1874), .b(n1873), .O(n1875));
  nand2 g1812(.a(n1875), .b(n1872), .O(n1876));
  nand2 g1813(.a(b15 ), .b(a8 ), .O(n1877));
  nand2 g1814(.a(b14 ), .b(a9 ), .O(n1878));
  inv1  g1815(.a(n1878), .O(n1879));
  nand2 g1816(.a(b13 ), .b(a10 ), .O(n1880));
  inv1  g1817(.a(n1880), .O(n1881));
  nand2 g1818(.a(b12 ), .b(a11 ), .O(n1882));
  inv1  g1819(.a(n1882), .O(n1883));
  nand2 g1820(.a(b11 ), .b(a12 ), .O(n1884));
  inv1  g1821(.a(n1884), .O(n1885));
  nand2 g1822(.a(b10 ), .b(a13 ), .O(n1886));
  inv1  g1823(.a(n1886), .O(n1887));
  nand2 g1824(.a(b9 ), .b(a14 ), .O(n1888));
  nand2 g1825(.a(b8 ), .b(a15 ), .O(n1889));
  xnor2 g1826(.a(n1889), .b(n1888), .O(n1890));
  inv1  g1827(.a(n1797), .O(n1891));
  nand2 g1828(.a(n1805), .b(n1891), .O(n1892));
  inv1  g1829(.a(n1796), .O(n1893));
  nand2 g1830(.a(n1805), .b(n1893), .O(n1894));
  nand2 g1831(.a(n1891), .b(n1893), .O(n1895));
  and2  g1832(.a(n1895), .b(n1894), .O(n1896));
  nand2 g1833(.a(n1896), .b(n1892), .O(n1897));
  xor2  g1834(.a(n1897), .b(n1890), .O(n1898));
  xor2  g1835(.a(n1898), .b(n1887), .O(n1899));
  inv1  g1836(.a(n1806), .O(n1900));
  nand2 g1837(.a(n1813), .b(n1900), .O(n1901));
  nand2 g1838(.a(n1813), .b(n1795), .O(n1902));
  nand2 g1839(.a(n1900), .b(n1795), .O(n1903));
  and2  g1840(.a(n1903), .b(n1902), .O(n1904));
  nand2 g1841(.a(n1904), .b(n1901), .O(n1905));
  xor2  g1842(.a(n1905), .b(n1899), .O(n1906));
  xor2  g1843(.a(n1906), .b(n1885), .O(n1907));
  inv1  g1844(.a(n1814), .O(n1908));
  nand2 g1845(.a(n1821), .b(n1908), .O(n1909));
  nand2 g1846(.a(n1821), .b(n1793), .O(n1910));
  nand2 g1847(.a(n1908), .b(n1793), .O(n1911));
  and2  g1848(.a(n1911), .b(n1910), .O(n1912));
  nand2 g1849(.a(n1912), .b(n1909), .O(n1913));
  xor2  g1850(.a(n1913), .b(n1907), .O(n1914));
  xor2  g1851(.a(n1914), .b(n1883), .O(n1915));
  inv1  g1852(.a(n1822), .O(n1916));
  nand2 g1853(.a(n1829), .b(n1916), .O(n1917));
  nand2 g1854(.a(n1829), .b(n1791), .O(n1918));
  nand2 g1855(.a(n1916), .b(n1791), .O(n1919));
  and2  g1856(.a(n1919), .b(n1918), .O(n1920));
  nand2 g1857(.a(n1920), .b(n1917), .O(n1921));
  xor2  g1858(.a(n1921), .b(n1915), .O(n1922));
  xor2  g1859(.a(n1922), .b(n1881), .O(n1923));
  inv1  g1860(.a(n1830), .O(n1924));
  nand2 g1861(.a(n1837), .b(n1924), .O(n1925));
  nand2 g1862(.a(n1837), .b(n1789), .O(n1926));
  nand2 g1863(.a(n1924), .b(n1789), .O(n1927));
  and2  g1864(.a(n1927), .b(n1926), .O(n1928));
  nand2 g1865(.a(n1928), .b(n1925), .O(n1929));
  xor2  g1866(.a(n1929), .b(n1923), .O(n1930));
  xor2  g1867(.a(n1930), .b(n1879), .O(n1931));
  inv1  g1868(.a(n1838), .O(n1932));
  nand2 g1869(.a(n1845), .b(n1932), .O(n1933));
  nand2 g1870(.a(n1845), .b(n1787), .O(n1934));
  nand2 g1871(.a(n1932), .b(n1787), .O(n1935));
  and2  g1872(.a(n1935), .b(n1934), .O(n1936));
  nand2 g1873(.a(n1936), .b(n1933), .O(n1937));
  xor2  g1874(.a(n1937), .b(n1931), .O(n1938));
  xor2  g1875(.a(n1938), .b(n1877), .O(n1939));
  inv1  g1876(.a(n1846), .O(n1940));
  nand2 g1877(.a(n1853), .b(n1940), .O(n1941));
  nand2 g1878(.a(n1853), .b(n1785), .O(n1942));
  nand2 g1879(.a(n1940), .b(n1785), .O(n1943));
  and2  g1880(.a(n1943), .b(n1942), .O(n1944));
  nand2 g1881(.a(n1944), .b(n1941), .O(n1945));
  xor2  g1882(.a(n1945), .b(n1939), .O(n1946));
  xor2  g1883(.a(n1946), .b(n1876), .O(n1947));
  inv1  g1884(.a(n1854), .O(n1948));
  nand2 g1885(.a(n1861), .b(n1948), .O(n1949));
  inv1  g1886(.a(n1783), .O(n1950));
  nand2 g1887(.a(n1861), .b(n1950), .O(n1951));
  nand2 g1888(.a(n1948), .b(n1950), .O(n1952));
  and2  g1889(.a(n1952), .b(n1951), .O(n1953));
  nand2 g1890(.a(n1953), .b(n1949), .O(n1954));
  xor2  g1891(.a(n1954), .b(n1947), .O(z23 ));
  nand2 g1892(.a(n1954), .b(n1876), .O(n1956));
  nand2 g1893(.a(n1954), .b(n1946), .O(n1957));
  nand2 g1894(.a(n1946), .b(n1876), .O(n1958));
  and2  g1895(.a(n1958), .b(n1957), .O(n1959));
  nand2 g1896(.a(n1959), .b(n1956), .O(n1960));
  nand2 g1897(.a(b15 ), .b(a9 ), .O(n1961));
  nand2 g1898(.a(b14 ), .b(a10 ), .O(n1962));
  inv1  g1899(.a(n1962), .O(n1963));
  nand2 g1900(.a(b13 ), .b(a11 ), .O(n1964));
  inv1  g1901(.a(n1964), .O(n1965));
  nand2 g1902(.a(b12 ), .b(a12 ), .O(n1966));
  inv1  g1903(.a(n1966), .O(n1967));
  nand2 g1904(.a(b11 ), .b(a13 ), .O(n1968));
  inv1  g1905(.a(n1968), .O(n1969));
  nand2 g1906(.a(b10 ), .b(a14 ), .O(n1970));
  nand2 g1907(.a(b9 ), .b(a15 ), .O(n1971));
  xnor2 g1908(.a(n1971), .b(n1970), .O(n1972));
  inv1  g1909(.a(n1889), .O(n1973));
  nand2 g1910(.a(n1897), .b(n1973), .O(n1974));
  inv1  g1911(.a(n1888), .O(n1975));
  nand2 g1912(.a(n1897), .b(n1975), .O(n1976));
  nand2 g1913(.a(n1973), .b(n1975), .O(n1977));
  and2  g1914(.a(n1977), .b(n1976), .O(n1978));
  nand2 g1915(.a(n1978), .b(n1974), .O(n1979));
  xor2  g1916(.a(n1979), .b(n1972), .O(n1980));
  xor2  g1917(.a(n1980), .b(n1969), .O(n1981));
  inv1  g1918(.a(n1898), .O(n1982));
  nand2 g1919(.a(n1905), .b(n1982), .O(n1983));
  nand2 g1920(.a(n1905), .b(n1887), .O(n1984));
  nand2 g1921(.a(n1982), .b(n1887), .O(n1985));
  and2  g1922(.a(n1985), .b(n1984), .O(n1986));
  nand2 g1923(.a(n1986), .b(n1983), .O(n1987));
  xor2  g1924(.a(n1987), .b(n1981), .O(n1988));
  xor2  g1925(.a(n1988), .b(n1967), .O(n1989));
  inv1  g1926(.a(n1906), .O(n1990));
  nand2 g1927(.a(n1913), .b(n1990), .O(n1991));
  nand2 g1928(.a(n1913), .b(n1885), .O(n1992));
  nand2 g1929(.a(n1990), .b(n1885), .O(n1993));
  and2  g1930(.a(n1993), .b(n1992), .O(n1994));
  nand2 g1931(.a(n1994), .b(n1991), .O(n1995));
  xor2  g1932(.a(n1995), .b(n1989), .O(n1996));
  xor2  g1933(.a(n1996), .b(n1965), .O(n1997));
  inv1  g1934(.a(n1914), .O(n1998));
  nand2 g1935(.a(n1921), .b(n1998), .O(n1999));
  nand2 g1936(.a(n1921), .b(n1883), .O(n2000));
  nand2 g1937(.a(n1998), .b(n1883), .O(n2001));
  and2  g1938(.a(n2001), .b(n2000), .O(n2002));
  nand2 g1939(.a(n2002), .b(n1999), .O(n2003));
  xor2  g1940(.a(n2003), .b(n1997), .O(n2004));
  xor2  g1941(.a(n2004), .b(n1963), .O(n2005));
  inv1  g1942(.a(n1922), .O(n2006));
  nand2 g1943(.a(n1929), .b(n2006), .O(n2007));
  nand2 g1944(.a(n1929), .b(n1881), .O(n2008));
  nand2 g1945(.a(n2006), .b(n1881), .O(n2009));
  and2  g1946(.a(n2009), .b(n2008), .O(n2010));
  nand2 g1947(.a(n2010), .b(n2007), .O(n2011));
  xor2  g1948(.a(n2011), .b(n2005), .O(n2012));
  xor2  g1949(.a(n2012), .b(n1961), .O(n2013));
  inv1  g1950(.a(n1930), .O(n2014));
  nand2 g1951(.a(n1937), .b(n2014), .O(n2015));
  nand2 g1952(.a(n1937), .b(n1879), .O(n2016));
  nand2 g1953(.a(n2014), .b(n1879), .O(n2017));
  and2  g1954(.a(n2017), .b(n2016), .O(n2018));
  nand2 g1955(.a(n2018), .b(n2015), .O(n2019));
  xor2  g1956(.a(n2019), .b(n2013), .O(n2020));
  xor2  g1957(.a(n2020), .b(n1960), .O(n2021));
  inv1  g1958(.a(n1938), .O(n2022));
  nand2 g1959(.a(n1945), .b(n2022), .O(n2023));
  inv1  g1960(.a(n1877), .O(n2024));
  nand2 g1961(.a(n1945), .b(n2024), .O(n2025));
  nand2 g1962(.a(n2022), .b(n2024), .O(n2026));
  and2  g1963(.a(n2026), .b(n2025), .O(n2027));
  nand2 g1964(.a(n2027), .b(n2023), .O(n2028));
  xor2  g1965(.a(n2028), .b(n2021), .O(z24 ));
  nand2 g1966(.a(n2028), .b(n1960), .O(n2030));
  nand2 g1967(.a(n2028), .b(n2020), .O(n2031));
  nand2 g1968(.a(n2020), .b(n1960), .O(n2032));
  and2  g1969(.a(n2032), .b(n2031), .O(n2033));
  nand2 g1970(.a(n2033), .b(n2030), .O(n2034));
  nand2 g1971(.a(b15 ), .b(a10 ), .O(n2035));
  nand2 g1972(.a(b14 ), .b(a11 ), .O(n2036));
  inv1  g1973(.a(n2036), .O(n2037));
  nand2 g1974(.a(b13 ), .b(a12 ), .O(n2038));
  inv1  g1975(.a(n2038), .O(n2039));
  nand2 g1976(.a(b12 ), .b(a13 ), .O(n2040));
  inv1  g1977(.a(n2040), .O(n2041));
  nand2 g1978(.a(b11 ), .b(a14 ), .O(n2042));
  nand2 g1979(.a(b10 ), .b(a15 ), .O(n2043));
  xnor2 g1980(.a(n2043), .b(n2042), .O(n2044));
  inv1  g1981(.a(n1971), .O(n2045));
  nand2 g1982(.a(n1979), .b(n2045), .O(n2046));
  inv1  g1983(.a(n1970), .O(n2047));
  nand2 g1984(.a(n1979), .b(n2047), .O(n2048));
  nand2 g1985(.a(n2045), .b(n2047), .O(n2049));
  and2  g1986(.a(n2049), .b(n2048), .O(n2050));
  nand2 g1987(.a(n2050), .b(n2046), .O(n2051));
  xor2  g1988(.a(n2051), .b(n2044), .O(n2052));
  xor2  g1989(.a(n2052), .b(n2041), .O(n2053));
  inv1  g1990(.a(n1980), .O(n2054));
  nand2 g1991(.a(n1987), .b(n2054), .O(n2055));
  nand2 g1992(.a(n1987), .b(n1969), .O(n2056));
  nand2 g1993(.a(n2054), .b(n1969), .O(n2057));
  and2  g1994(.a(n2057), .b(n2056), .O(n2058));
  nand2 g1995(.a(n2058), .b(n2055), .O(n2059));
  xor2  g1996(.a(n2059), .b(n2053), .O(n2060));
  xor2  g1997(.a(n2060), .b(n2039), .O(n2061));
  inv1  g1998(.a(n1988), .O(n2062));
  nand2 g1999(.a(n1995), .b(n2062), .O(n2063));
  nand2 g2000(.a(n1995), .b(n1967), .O(n2064));
  nand2 g2001(.a(n2062), .b(n1967), .O(n2065));
  and2  g2002(.a(n2065), .b(n2064), .O(n2066));
  nand2 g2003(.a(n2066), .b(n2063), .O(n2067));
  xor2  g2004(.a(n2067), .b(n2061), .O(n2068));
  xor2  g2005(.a(n2068), .b(n2037), .O(n2069));
  inv1  g2006(.a(n1996), .O(n2070));
  nand2 g2007(.a(n2003), .b(n2070), .O(n2071));
  nand2 g2008(.a(n2003), .b(n1965), .O(n2072));
  nand2 g2009(.a(n2070), .b(n1965), .O(n2073));
  and2  g2010(.a(n2073), .b(n2072), .O(n2074));
  nand2 g2011(.a(n2074), .b(n2071), .O(n2075));
  xor2  g2012(.a(n2075), .b(n2069), .O(n2076));
  xor2  g2013(.a(n2076), .b(n2035), .O(n2077));
  inv1  g2014(.a(n2004), .O(n2078));
  nand2 g2015(.a(n2011), .b(n2078), .O(n2079));
  nand2 g2016(.a(n2011), .b(n1963), .O(n2080));
  nand2 g2017(.a(n2078), .b(n1963), .O(n2081));
  and2  g2018(.a(n2081), .b(n2080), .O(n2082));
  nand2 g2019(.a(n2082), .b(n2079), .O(n2083));
  xor2  g2020(.a(n2083), .b(n2077), .O(n2084));
  xor2  g2021(.a(n2084), .b(n2034), .O(n2085));
  inv1  g2022(.a(n2012), .O(n2086));
  nand2 g2023(.a(n2019), .b(n2086), .O(n2087));
  inv1  g2024(.a(n1961), .O(n2088));
  nand2 g2025(.a(n2019), .b(n2088), .O(n2089));
  nand2 g2026(.a(n2086), .b(n2088), .O(n2090));
  and2  g2027(.a(n2090), .b(n2089), .O(n2091));
  nand2 g2028(.a(n2091), .b(n2087), .O(n2092));
  xor2  g2029(.a(n2092), .b(n2085), .O(z25 ));
  nand2 g2030(.a(n2092), .b(n2034), .O(n2094));
  nand2 g2031(.a(n2092), .b(n2084), .O(n2095));
  nand2 g2032(.a(n2084), .b(n2034), .O(n2096));
  and2  g2033(.a(n2096), .b(n2095), .O(n2097));
  nand2 g2034(.a(n2097), .b(n2094), .O(n2098));
  nand2 g2035(.a(b15 ), .b(a11 ), .O(n2099));
  nand2 g2036(.a(b14 ), .b(a12 ), .O(n2100));
  inv1  g2037(.a(n2100), .O(n2101));
  nand2 g2038(.a(b13 ), .b(a13 ), .O(n2102));
  inv1  g2039(.a(n2102), .O(n2103));
  nand2 g2040(.a(b12 ), .b(a14 ), .O(n2104));
  nand2 g2041(.a(b11 ), .b(a15 ), .O(n2105));
  xnor2 g2042(.a(n2105), .b(n2104), .O(n2106));
  inv1  g2043(.a(n2043), .O(n2107));
  nand2 g2044(.a(n2051), .b(n2107), .O(n2108));
  inv1  g2045(.a(n2042), .O(n2109));
  nand2 g2046(.a(n2051), .b(n2109), .O(n2110));
  nand2 g2047(.a(n2107), .b(n2109), .O(n2111));
  and2  g2048(.a(n2111), .b(n2110), .O(n2112));
  nand2 g2049(.a(n2112), .b(n2108), .O(n2113));
  xor2  g2050(.a(n2113), .b(n2106), .O(n2114));
  xor2  g2051(.a(n2114), .b(n2103), .O(n2115));
  inv1  g2052(.a(n2052), .O(n2116));
  nand2 g2053(.a(n2059), .b(n2116), .O(n2117));
  nand2 g2054(.a(n2059), .b(n2041), .O(n2118));
  nand2 g2055(.a(n2116), .b(n2041), .O(n2119));
  and2  g2056(.a(n2119), .b(n2118), .O(n2120));
  nand2 g2057(.a(n2120), .b(n2117), .O(n2121));
  xor2  g2058(.a(n2121), .b(n2115), .O(n2122));
  xor2  g2059(.a(n2122), .b(n2101), .O(n2123));
  inv1  g2060(.a(n2060), .O(n2124));
  nand2 g2061(.a(n2067), .b(n2124), .O(n2125));
  nand2 g2062(.a(n2067), .b(n2039), .O(n2126));
  nand2 g2063(.a(n2124), .b(n2039), .O(n2127));
  and2  g2064(.a(n2127), .b(n2126), .O(n2128));
  nand2 g2065(.a(n2128), .b(n2125), .O(n2129));
  xor2  g2066(.a(n2129), .b(n2123), .O(n2130));
  xor2  g2067(.a(n2130), .b(n2099), .O(n2131));
  inv1  g2068(.a(n2068), .O(n2132));
  nand2 g2069(.a(n2075), .b(n2132), .O(n2133));
  nand2 g2070(.a(n2075), .b(n2037), .O(n2134));
  nand2 g2071(.a(n2132), .b(n2037), .O(n2135));
  and2  g2072(.a(n2135), .b(n2134), .O(n2136));
  nand2 g2073(.a(n2136), .b(n2133), .O(n2137));
  xor2  g2074(.a(n2137), .b(n2131), .O(n2138));
  xor2  g2075(.a(n2138), .b(n2098), .O(n2139));
  inv1  g2076(.a(n2076), .O(n2140));
  nand2 g2077(.a(n2083), .b(n2140), .O(n2141));
  inv1  g2078(.a(n2035), .O(n2142));
  nand2 g2079(.a(n2083), .b(n2142), .O(n2143));
  nand2 g2080(.a(n2140), .b(n2142), .O(n2144));
  and2  g2081(.a(n2144), .b(n2143), .O(n2145));
  nand2 g2082(.a(n2145), .b(n2141), .O(n2146));
  xor2  g2083(.a(n2146), .b(n2139), .O(z26 ));
  nand2 g2084(.a(n2146), .b(n2098), .O(n2148));
  nand2 g2085(.a(n2146), .b(n2138), .O(n2149));
  nand2 g2086(.a(n2138), .b(n2098), .O(n2150));
  and2  g2087(.a(n2150), .b(n2149), .O(n2151));
  nand2 g2088(.a(n2151), .b(n2148), .O(n2152));
  nand2 g2089(.a(b15 ), .b(a12 ), .O(n2153));
  nand2 g2090(.a(b14 ), .b(a13 ), .O(n2154));
  inv1  g2091(.a(n2154), .O(n2155));
  nand2 g2092(.a(b13 ), .b(a14 ), .O(n2156));
  nand2 g2093(.a(b12 ), .b(a15 ), .O(n2157));
  xnor2 g2094(.a(n2157), .b(n2156), .O(n2158));
  inv1  g2095(.a(n2105), .O(n2159));
  nand2 g2096(.a(n2113), .b(n2159), .O(n2160));
  inv1  g2097(.a(n2104), .O(n2161));
  nand2 g2098(.a(n2113), .b(n2161), .O(n2162));
  nand2 g2099(.a(n2159), .b(n2161), .O(n2163));
  and2  g2100(.a(n2163), .b(n2162), .O(n2164));
  nand2 g2101(.a(n2164), .b(n2160), .O(n2165));
  xor2  g2102(.a(n2165), .b(n2158), .O(n2166));
  xor2  g2103(.a(n2166), .b(n2155), .O(n2167));
  inv1  g2104(.a(n2114), .O(n2168));
  nand2 g2105(.a(n2121), .b(n2168), .O(n2169));
  nand2 g2106(.a(n2121), .b(n2103), .O(n2170));
  nand2 g2107(.a(n2168), .b(n2103), .O(n2171));
  and2  g2108(.a(n2171), .b(n2170), .O(n2172));
  nand2 g2109(.a(n2172), .b(n2169), .O(n2173));
  xor2  g2110(.a(n2173), .b(n2167), .O(n2174));
  xor2  g2111(.a(n2174), .b(n2153), .O(n2175));
  inv1  g2112(.a(n2122), .O(n2176));
  nand2 g2113(.a(n2129), .b(n2176), .O(n2177));
  nand2 g2114(.a(n2129), .b(n2101), .O(n2178));
  nand2 g2115(.a(n2176), .b(n2101), .O(n2179));
  and2  g2116(.a(n2179), .b(n2178), .O(n2180));
  nand2 g2117(.a(n2180), .b(n2177), .O(n2181));
  xor2  g2118(.a(n2181), .b(n2175), .O(n2182));
  xor2  g2119(.a(n2182), .b(n2152), .O(n2183));
  inv1  g2120(.a(n2130), .O(n2184));
  nand2 g2121(.a(n2137), .b(n2184), .O(n2185));
  inv1  g2122(.a(n2099), .O(n2186));
  nand2 g2123(.a(n2137), .b(n2186), .O(n2187));
  nand2 g2124(.a(n2184), .b(n2186), .O(n2188));
  and2  g2125(.a(n2188), .b(n2187), .O(n2189));
  nand2 g2126(.a(n2189), .b(n2185), .O(n2190));
  xor2  g2127(.a(n2190), .b(n2183), .O(z27 ));
  nand2 g2128(.a(n2190), .b(n2152), .O(n2192));
  nand2 g2129(.a(n2190), .b(n2182), .O(n2193));
  nand2 g2130(.a(n2182), .b(n2152), .O(n2194));
  and2  g2131(.a(n2194), .b(n2193), .O(n2195));
  nand2 g2132(.a(n2195), .b(n2192), .O(n2196));
  nand2 g2133(.a(b15 ), .b(a13 ), .O(n2197));
  nand2 g2134(.a(b14 ), .b(a14 ), .O(n2198));
  nand2 g2135(.a(b13 ), .b(a15 ), .O(n2199));
  xnor2 g2136(.a(n2199), .b(n2198), .O(n2200));
  inv1  g2137(.a(n2157), .O(n2201));
  nand2 g2138(.a(n2165), .b(n2201), .O(n2202));
  inv1  g2139(.a(n2156), .O(n2203));
  nand2 g2140(.a(n2165), .b(n2203), .O(n2204));
  nand2 g2141(.a(n2201), .b(n2203), .O(n2205));
  and2  g2142(.a(n2205), .b(n2204), .O(n2206));
  nand2 g2143(.a(n2206), .b(n2202), .O(n2207));
  xor2  g2144(.a(n2207), .b(n2200), .O(n2208));
  xor2  g2145(.a(n2208), .b(n2197), .O(n2209));
  inv1  g2146(.a(n2166), .O(n2210));
  nand2 g2147(.a(n2173), .b(n2210), .O(n2211));
  nand2 g2148(.a(n2173), .b(n2155), .O(n2212));
  nand2 g2149(.a(n2210), .b(n2155), .O(n2213));
  and2  g2150(.a(n2213), .b(n2212), .O(n2214));
  nand2 g2151(.a(n2214), .b(n2211), .O(n2215));
  xor2  g2152(.a(n2215), .b(n2209), .O(n2216));
  xor2  g2153(.a(n2216), .b(n2196), .O(n2217));
  inv1  g2154(.a(n2174), .O(n2218));
  nand2 g2155(.a(n2181), .b(n2218), .O(n2219));
  inv1  g2156(.a(n2153), .O(n2220));
  nand2 g2157(.a(n2181), .b(n2220), .O(n2221));
  nand2 g2158(.a(n2218), .b(n2220), .O(n2222));
  and2  g2159(.a(n2222), .b(n2221), .O(n2223));
  nand2 g2160(.a(n2223), .b(n2219), .O(n2224));
  xor2  g2161(.a(n2224), .b(n2217), .O(z28 ));
  nand2 g2162(.a(n2224), .b(n2196), .O(n2226));
  nand2 g2163(.a(n2224), .b(n2216), .O(n2227));
  nand2 g2164(.a(n2216), .b(n2196), .O(n2228));
  and2  g2165(.a(n2228), .b(n2227), .O(n2229));
  nand2 g2166(.a(n2229), .b(n2226), .O(n2230));
  nand2 g2167(.a(b15 ), .b(a14 ), .O(n2231));
  nand2 g2168(.a(b14 ), .b(a15 ), .O(n2232));
  xor2  g2169(.a(n2232), .b(n2231), .O(n2233));
  inv1  g2170(.a(n2199), .O(n2234));
  nand2 g2171(.a(n2207), .b(n2234), .O(n2235));
  inv1  g2172(.a(n2198), .O(n2236));
  nand2 g2173(.a(n2207), .b(n2236), .O(n2237));
  nand2 g2174(.a(n2234), .b(n2236), .O(n2238));
  and2  g2175(.a(n2238), .b(n2237), .O(n2239));
  nand2 g2176(.a(n2239), .b(n2235), .O(n2240));
  xor2  g2177(.a(n2240), .b(n2233), .O(n2241));
  xor2  g2178(.a(n2241), .b(n2230), .O(n2242));
  inv1  g2179(.a(n2208), .O(n2243));
  nand2 g2180(.a(n2215), .b(n2243), .O(n2244));
  inv1  g2181(.a(n2197), .O(n2245));
  nand2 g2182(.a(n2215), .b(n2245), .O(n2246));
  nand2 g2183(.a(n2243), .b(n2245), .O(n2247));
  and2  g2184(.a(n2247), .b(n2246), .O(n2248));
  nand2 g2185(.a(n2248), .b(n2244), .O(n2249));
  xor2  g2186(.a(n2249), .b(n2242), .O(z29 ));
  nand2 g2187(.a(n2249), .b(n2230), .O(n2251));
  nand2 g2188(.a(n2249), .b(n2241), .O(n2252));
  nand2 g2189(.a(n2241), .b(n2230), .O(n2253));
  and2  g2190(.a(n2253), .b(n2252), .O(n2254));
  nand2 g2191(.a(n2254), .b(n2251), .O(n2255));
  and2  g2192(.a(b15 ), .b(a15 ), .O(n2256));
  xor2  g2193(.a(n2256), .b(n2255), .O(n2257));
  inv1  g2194(.a(n2232), .O(n2258));
  nand2 g2195(.a(n2240), .b(n2258), .O(n2259));
  inv1  g2196(.a(n2231), .O(n2260));
  nand2 g2197(.a(n2240), .b(n2260), .O(n2261));
  nand2 g2198(.a(n2258), .b(n2260), .O(n2262));
  and2  g2199(.a(n2262), .b(n2261), .O(n2263));
  nand2 g2200(.a(n2263), .b(n2259), .O(n2264));
  xor2  g2201(.a(n2264), .b(n2257), .O(z30 ));
  nand2 g2202(.a(n2264), .b(n2255), .O(n2266));
  nand2 g2203(.a(n2264), .b(n2256), .O(n2267));
  nand2 g2204(.a(n2256), .b(n2255), .O(n2268));
  and2  g2205(.a(n2268), .b(n2267), .O(n2269));
  nand2 g2206(.a(n2269), .b(n2266), .O(z31 ));
endmodule


